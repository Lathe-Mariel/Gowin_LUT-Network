`timescale 1ns / 1ps



module MnistLutSimple
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire                  reset,
            input  wire                  clk,
            input  wire                  cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [      784-1:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [       10-1:0]  out_data,
            output wire                  out_valid
        );
    
    
    wire  [USER_BITS-1:0]  layer0_user;
    wire  [     1024-1:0]  layer0_data;
    wire                   layer0_valid;
    
    MnistLutSimple_sub0
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub0
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (in_user),
                .in_data    (in_data),
                .in_valid   (in_valid),
                
                .out_user   (layer0_user),
                .out_data   (layer0_data),
                .out_valid  (layer0_valid)
             );
    
    wire  [USER_BITS-1:0]  layer1_user;
    wire  [      512-1:0]  layer1_data;
    wire                   layer1_valid;
    
    MnistLutSimple_sub1
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub1
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer0_user),
                .in_data    (layer0_data),
                .in_valid   (layer0_valid),
                
                .out_user   (layer1_user),
                .out_data   (layer1_data),
                .out_valid  (layer1_valid)
             );
    
    wire  [USER_BITS-1:0]  layer2_user;
    wire  [      640-1:0]  layer2_data;
    wire                   layer2_valid;
    
    MnistLutSimple_sub2
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub2
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer1_user),
                .in_data    (layer1_data),
                .in_valid   (layer1_valid),
                
                .out_user   (layer2_user),
                .out_data   (layer2_data),
                .out_valid  (layer2_valid)
             );
    
    wire  [USER_BITS-1:0]  layer3_user;
    wire  [      640-1:0]  layer3_data;
    wire                   layer3_valid;
    
    MnistLutSimple_sub3
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub3
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer2_user),
                .in_data    (layer2_data),
                .in_valid   (layer2_valid),
                
                .out_user   (layer3_user),
                .out_data   (layer3_data),
                .out_valid  (layer3_valid)
             );
    
    wire  [USER_BITS-1:0]  layer4_user;
    wire  [      640-1:0]  layer4_data;
    wire                   layer4_valid;
    
    MnistLutSimple_sub4
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub4
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer3_user),
                .in_data    (layer3_data),
                .in_valid   (layer3_valid),
                
                .out_user   (layer4_user),
                .out_data   (layer4_data),
                .out_valid  (layer4_valid)
             );
    
    wire  [USER_BITS-1:0]  layer5_user;
    wire  [      640-1:0]  layer5_data;
    wire                   layer5_valid;
    
    MnistLutSimple_sub5
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub5
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer4_user),
                .in_data    (layer4_data),
                .in_valid   (layer4_valid),
                
                .out_user   (layer5_user),
                .out_data   (layer5_data),
                .out_valid  (layer5_valid)
             );
    
    wire  [USER_BITS-1:0]  layer6_user;
    wire  [      160-1:0]  layer6_data;
    wire                   layer6_valid;
    
    MnistLutSimple_sub6
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub6
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer5_user),
                .in_data    (layer5_data),
                .in_valid   (layer5_valid),
                
                .out_user   (layer6_user),
                .out_data   (layer6_data),
                .out_valid  (layer6_valid)
             );
    
    wire  [USER_BITS-1:0]  layer7_user;
    wire  [       40-1:0]  layer7_data;
    wire                   layer7_valid;
    
    MnistLutSimple_sub7
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub7
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer6_user),
                .in_data    (layer6_data),
                .in_valid   (layer6_valid),
                
                .out_user   (layer7_user),
                .out_data   (layer7_data),
                .out_valid  (layer7_valid)
             );
    
    wire  [USER_BITS-1:0]  layer8_user;
    wire  [       10-1:0]  layer8_data;
    wire                   layer8_valid;
    
    MnistLutSimple_sub8
            #(
                .USER_WIDTH (USER_WIDTH),
                .USE_REG    (USE_REG),
                .INIT_REG   (INIT_REG),
                .DEVICE     (DEVICE)
            )
        i_MnistLutSimple_sub8
            (
                .reset      (reset),
                .clk        (clk),
                .cke        (cke),
                
                .in_user    (layer7_user),
                .in_data    (layer7_data),
                .in_valid   (layer7_valid),
                
                .out_user   (layer8_user),
                .out_data   (layer8_data),
                .out_valid  (layer8_valid)
             );
    
    assign out_data  = layer8_data;
    assign out_user  = layer8_user;
    assign out_valid = layer8_valid;
    
endmodule




module MnistLutSimple_sub0
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        783:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [       1023:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub0_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub0_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub0_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [783:0]  in_data,
            output wire [1023:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1111101011101111;
    wire [3:0] lut_0_select = {
                             in_data[459],
                             in_data[432],
                             in_data[227],
                             in_data[285]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b1111111011111110;
    wire [3:0] lut_1_select = {
                             in_data[4],
                             in_data[246],
                             in_data[502],
                             in_data[774]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b0000000001011001;
    wire [3:0] lut_2_select = {
                             in_data[638],
                             in_data[287],
                             in_data[633],
                             in_data[148]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1111111111111110;
    wire [3:0] lut_3_select = {
                             in_data[507],
                             in_data[175],
                             in_data[679],
                             in_data[590]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b0101010100000101;
    wire [3:0] lut_4_select = {
                             in_data[413],
                             in_data[153],
                             in_data[196],
                             in_data[123]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1111111111011100;
    wire [3:0] lut_5_select = {
                             in_data[99],
                             in_data[212],
                             in_data[608],
                             in_data[105]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b0100010001000100;
    wire [3:0] lut_6_select = {
                             in_data[71],
                             in_data[775],
                             in_data[653],
                             in_data[735]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b0000111100001111;
    wire [3:0] lut_7_select = {
                             in_data[357],
                             in_data[659],
                             in_data[419],
                             in_data[699]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1111111111111100;
    wire [3:0] lut_8_select = {
                             in_data[606],
                             in_data[247],
                             in_data[472],
                             in_data[19]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b0010000011111111;
    wire [3:0] lut_9_select = {
                             in_data[211],
                             in_data[586],
                             in_data[163],
                             in_data[769]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b1111111100001010;
    wire [3:0] lut_10_select = {
                             in_data[569],
                             in_data[381],
                             in_data[761],
                             in_data[647]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b0011001100110000;
    wire [3:0] lut_11_select = {
                             in_data[282],
                             in_data[438],
                             in_data[360],
                             in_data[113]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b1111110011111101;
    wire [3:0] lut_12_select = {
                             in_data[727],
                             in_data[451],
                             in_data[744],
                             in_data[585]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0000000011111111;
    wire [3:0] lut_13_select = {
                             in_data[155],
                             in_data[293],
                             in_data[573],
                             in_data[674]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0111001101110011;
    wire [3:0] lut_14_select = {
                             in_data[760],
                             in_data[146],
                             in_data[292],
                             in_data[192]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1111110111110100;
    wire [3:0] lut_15_select = {
                             in_data[92],
                             in_data[388],
                             in_data[603],
                             in_data[430]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b1111111110110000;
    wire [3:0] lut_16_select = {
                             in_data[93],
                             in_data[575],
                             in_data[464],
                             in_data[232]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b0000111100001111;
    wire [3:0] lut_17_select = {
                             in_data[520],
                             in_data[300],
                             in_data[107],
                             in_data[504]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0101010101010101;
    wire [3:0] lut_18_select = {
                             in_data[242],
                             in_data[161],
                             in_data[533],
                             in_data[324]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b1111111111110000;
    wire [3:0] lut_19_select = {
                             in_data[129],
                             in_data[594],
                             in_data[330],
                             in_data[114]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0000010001000100;
    wire [3:0] lut_20_select = {
                             in_data[144],
                             in_data[637],
                             in_data[684],
                             in_data[183]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b0000000100110101;
    wire [3:0] lut_21_select = {
                             in_data[185],
                             in_data[191],
                             in_data[170],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b0000101100001011;
    wire [3:0] lut_22_select = {
                             in_data[778],
                             in_data[220],
                             in_data[371],
                             in_data[261]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b1111000011110110;
    wire [3:0] lut_23_select = {
                             in_data[409],
                             in_data[178],
                             in_data[686],
                             in_data[498]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1111011101010000;
    wire [3:0] lut_24_select = {
                             in_data[34],
                             in_data[122],
                             in_data[696],
                             in_data[776]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0000010001010101;
    wire [3:0] lut_25_select = {
                             in_data[296],
                             in_data[591],
                             in_data[598],
                             in_data[424]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b0000010100000101;
    wire [3:0] lut_26_select = {
                             in_data[313],
                             in_data[154],
                             in_data[530],
                             in_data[570]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1111111111111110;
    wire [3:0] lut_27_select = {
                             in_data[222],
                             in_data[609],
                             in_data[280],
                             in_data[66]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b1010111110101111;
    wire [3:0] lut_28_select = {
                             in_data[667],
                             in_data[494],
                             in_data[140],
                             in_data[69]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b1000101100001111;
    wire [3:0] lut_29_select = {
                             in_data[37],
                             in_data[180],
                             in_data[600],
                             in_data[532]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b1010000010100001;
    wire [3:0] lut_30_select = {
                             in_data[40],
                             in_data[514],
                             in_data[64],
                             in_data[453]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b0000101010101110;
    wire [3:0] lut_31_select = {
                             in_data[648],
                             in_data[230],
                             in_data[528],
                             in_data[455]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1111111100001111;
    wire [3:0] lut_32_select = {
                             in_data[583],
                             in_data[260],
                             in_data[560],
                             in_data[666]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b1100111111001111;
    wire [3:0] lut_33_select = {
                             in_data[24],
                             in_data[461],
                             in_data[68],
                             in_data[703]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1111111111111100;
    wire [3:0] lut_34_select = {
                             in_data[350],
                             in_data[307],
                             in_data[120],
                             in_data[20]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1111111111101110;
    wire [3:0] lut_35_select = {
                             in_data[554],
                             in_data[751],
                             in_data[595],
                             in_data[563]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b1101110100001000;
    wire [3:0] lut_36_select = {
                             in_data[431],
                             in_data[386],
                             in_data[354],
                             in_data[164]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0000000000110010;
    wire [3:0] lut_37_select = {
                             in_data[284],
                             in_data[643],
                             in_data[139],
                             in_data[26]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b0010001010101010;
    wire [3:0] lut_38_select = {
                             in_data[204],
                             in_data[725],
                             in_data[465],
                             in_data[210]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0100110011001101;
    wire [3:0] lut_39_select = {
                             in_data[397],
                             in_data[390],
                             in_data[97],
                             in_data[773]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b1111110011111100;
    wire [3:0] lut_40_select = {
                             in_data[753],
                             in_data[500],
                             in_data[104],
                             in_data[422]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b0000110100001111;
    wire [3:0] lut_41_select = {
                             in_data[645],
                             in_data[688],
                             in_data[538],
                             in_data[111]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b0100110101000101;
    wire [3:0] lut_42_select = {
                             in_data[336],
                             in_data[171],
                             in_data[395],
                             in_data[270]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0000000100000001;
    wire [3:0] lut_43_select = {
                             in_data[11],
                             in_data[711],
                             in_data[301],
                             in_data[394]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b1111101011111011;
    wire [3:0] lut_44_select = {
                             in_data[50],
                             in_data[478],
                             in_data[233],
                             in_data[709]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b0101010100000000;
    wire [3:0] lut_45_select = {
                             in_data[238],
                             in_data[671],
                             in_data[138],
                             in_data[486]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b1100010011000100;
    wire [3:0] lut_46_select = {
                             in_data[450],
                             in_data[434],
                             in_data[517],
                             in_data[546]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b0100010001000100;
    wire [3:0] lut_47_select = {
                             in_data[9],
                             in_data[1],
                             in_data[383],
                             in_data[278]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b0000001000000010;
    wire [3:0] lut_48_select = {
                             in_data[224],
                             in_data[249],
                             in_data[693],
                             in_data[739]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b0010101000101010;
    wire [3:0] lut_49_select = {
                             in_data[759],
                             in_data[721],
                             in_data[124],
                             in_data[541]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0011000011111111;
    wire [3:0] lut_50_select = {
                             in_data[518],
                             in_data[197],
                             in_data[471],
                             in_data[561]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b1000100011111111;
    wire [3:0] lut_51_select = {
                             in_data[240],
                             in_data[589],
                             in_data[635],
                             in_data[750]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1111111100010001;
    wire [3:0] lut_52_select = {
                             in_data[715],
                             in_data[30],
                             in_data[661],
                             in_data[339]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b0001000000110000;
    wire [3:0] lut_53_select = {
                             in_data[477],
                             in_data[147],
                             in_data[640],
                             in_data[62]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b0000000001010000;
    wire [3:0] lut_54_select = {
                             in_data[580],
                             in_data[346],
                             in_data[168],
                             in_data[203]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b1111111111111110;
    wire [3:0] lut_55_select = {
                             in_data[558],
                             in_data[226],
                             in_data[487],
                             in_data[488]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b1111000011110000;
    wire [3:0] lut_56_select = {
                             in_data[5],
                             in_data[298],
                             in_data[127],
                             in_data[476]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b1111111111110000;
    wire [3:0] lut_57_select = {
                             in_data[454],
                             in_data[315],
                             in_data[448],
                             in_data[27]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b0001000100000000;
    wire [3:0] lut_58_select = {
                             in_data[463],
                             in_data[65],
                             in_data[649],
                             in_data[255]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b1111111110101010;
    wire [3:0] lut_59_select = {
                             in_data[160],
                             in_data[45],
                             in_data[698],
                             in_data[539]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b0000010100000101;
    wire [3:0] lut_60_select = {
                             in_data[28],
                             in_data[391],
                             in_data[529],
                             in_data[762]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b0000001100000000;
    wire [3:0] lut_61_select = {
                             in_data[345],
                             in_data[581],
                             in_data[738],
                             in_data[481]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b0101010100000000;
    wire [3:0] lut_62_select = {
                             in_data[480],
                             in_data[425],
                             in_data[250],
                             in_data[396]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b1111000011111101;
    wire [3:0] lut_63_select = {
                             in_data[248],
                             in_data[708],
                             in_data[663],
                             in_data[700]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b0001000100010001;
    wire [3:0] lut_64_select = {
                             in_data[690],
                             in_data[88],
                             in_data[442],
                             in_data[439]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b0010000000000101;
    wire [3:0] lut_65_select = {
                             in_data[437],
                             in_data[95],
                             in_data[17],
                             in_data[382]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b1111111111111110;
    wire [3:0] lut_66_select = {
                             in_data[564],
                             in_data[179],
                             in_data[121],
                             in_data[510]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b1110111011101110;
    wire [3:0] lut_67_select = {
                             in_data[7],
                             in_data[59],
                             in_data[332],
                             in_data[374]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b1010000011111111;
    wire [3:0] lut_68_select = {
                             in_data[491],
                             in_data[402],
                             in_data[616],
                             in_data[676]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b0010000010110000;
    wire [3:0] lut_69_select = {
                             in_data[254],
                             in_data[209],
                             in_data[446],
                             in_data[239]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b0110011000000101;
    wire [3:0] lut_70_select = {
                             in_data[599],
                             in_data[256],
                             in_data[231],
                             in_data[547]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b1011111010101110;
    wire [3:0] lut_71_select = {
                             in_data[612],
                             in_data[152],
                             in_data[410],
                             in_data[710]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b0011000000110011;
    wire [3:0] lut_72_select = {
                             in_data[131],
                             in_data[143],
                             in_data[660],
                             in_data[726]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b1011101100000000;
    wire [3:0] lut_73_select = {
                             in_data[657],
                             in_data[13],
                             in_data[337],
                             in_data[662]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0000000011011101;
    wire [3:0] lut_74_select = {
                             in_data[400],
                             in_data[12],
                             in_data[605],
                             in_data[764]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b1111101011111010;
    wire [3:0] lut_75_select = {
                             in_data[23],
                             in_data[362],
                             in_data[162],
                             in_data[537]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0000110111001101;
    wire [3:0] lut_76_select = {
                             in_data[376],
                             in_data[94],
                             in_data[331],
                             in_data[492]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b0100010001001100;
    wire [3:0] lut_77_select = {
                             in_data[286],
                             in_data[683],
                             in_data[358],
                             in_data[257]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b0000000001010101;
    wire [3:0] lut_78_select = {
                             in_data[513],
                             in_data[697],
                             in_data[617],
                             in_data[565]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b1101110111111101;
    wire [3:0] lut_79_select = {
                             in_data[577],
                             in_data[694],
                             in_data[452],
                             in_data[630]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b0100010001000100;
    wire [3:0] lut_80_select = {
                             in_data[615],
                             in_data[87],
                             in_data[351],
                             in_data[678]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b1100110011111110;
    wire [3:0] lut_81_select = {
                             in_data[691],
                             in_data[550],
                             in_data[172],
                             in_data[493]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b0000000000010001;
    wire [3:0] lut_82_select = {
                             in_data[720],
                             in_data[108],
                             in_data[317],
                             in_data[717]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b0000101000000000;
    wire [3:0] lut_83_select = {
                             in_data[291],
                             in_data[258],
                             in_data[613],
                             in_data[320]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b0001000100000000;
    wire [3:0] lut_84_select = {
                             in_data[323],
                             in_data[749],
                             in_data[259],
                             in_data[289]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b1000111011101110;
    wire [3:0] lut_85_select = {
                             in_data[311],
                             in_data[629],
                             in_data[523],
                             in_data[457]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b1111111100001111;
    wire [3:0] lut_86_select = {
                             in_data[770],
                             in_data[496],
                             in_data[335],
                             in_data[333]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b1111110011111100;
    wire [3:0] lut_87_select = {
                             in_data[596],
                             in_data[375],
                             in_data[398],
                             in_data[754]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b1111111111111100;
    wire [3:0] lut_88_select = {
                             in_data[135],
                             in_data[253],
                             in_data[423],
                             in_data[475]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b1111111111111100;
    wire [3:0] lut_89_select = {
                             in_data[283],
                             in_data[117],
                             in_data[265],
                             in_data[706]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1111111110101110;
    wire [3:0] lut_90_select = {
                             in_data[126],
                             in_data[522],
                             in_data[729],
                             in_data[445]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b0000000001010000;
    wire [3:0] lut_91_select = {
                             in_data[200],
                             in_data[406],
                             in_data[194],
                             in_data[468]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1101110111011101;
    wire [3:0] lut_92_select = {
                             in_data[201],
                             in_data[695],
                             in_data[219],
                             in_data[404]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0000000000000011;
    wire [3:0] lut_93_select = {
                             in_data[96],
                             in_data[650],
                             in_data[15],
                             in_data[6]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b1010101000001101;
    wire [3:0] lut_94_select = {
                             in_data[150],
                             in_data[552],
                             in_data[625],
                             in_data[263]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b1111101011111111;
    wire [3:0] lut_95_select = {
                             in_data[85],
                             in_data[780],
                             in_data[783],
                             in_data[766]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1111000011110000;
    wire [3:0] lut_96_select = {
                             in_data[642],
                             in_data[319],
                             in_data[89],
                             in_data[288]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b0000000010110010;
    wire [3:0] lut_97_select = {
                             in_data[473],
                             in_data[444],
                             in_data[677],
                             in_data[628]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1010101011101110;
    wire [3:0] lut_98_select = {
                             in_data[262],
                             in_data[166],
                             in_data[495],
                             in_data[639]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b1111000011111100;
    wire [3:0] lut_99_select = {
                             in_data[752],
                             in_data[101],
                             in_data[379],
                             in_data[141]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1100110111001101;
    wire [3:0] lut_100_select = {
                             in_data[32],
                             in_data[571],
                             in_data[145],
                             in_data[49]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b0000010100000101;
    wire [3:0] lut_101_select = {
                             in_data[0],
                             in_data[470],
                             in_data[420],
                             in_data[733]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b1010111011111111;
    wire [3:0] lut_102_select = {
                             in_data[213],
                             in_data[393],
                             in_data[86],
                             in_data[142]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1010111100101111;
    wire [3:0] lut_103_select = {
                             in_data[77],
                             in_data[369],
                             in_data[556],
                             in_data[416]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b1111111111111110;
    wire [3:0] lut_104_select = {
                             in_data[622],
                             in_data[314],
                             in_data[719],
                             in_data[356]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1000111110101010;
    wire [3:0] lut_105_select = {
                             in_data[509],
                             in_data[190],
                             in_data[167],
                             in_data[544]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b0011001110110011;
    wire [3:0] lut_106_select = {
                             in_data[736],
                             in_data[748],
                             in_data[658],
                             in_data[427]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b0100010000110011;
    wire [3:0] lut_107_select = {
                             in_data[322],
                             in_data[728],
                             in_data[682],
                             in_data[159]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b1111111101001100;
    wire [3:0] lut_108_select = {
                             in_data[515],
                             in_data[574],
                             in_data[325],
                             in_data[519]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b1111110000111111;
    wire [3:0] lut_109_select = {
                             in_data[436],
                             in_data[125],
                             in_data[593],
                             in_data[29]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b1010111010101110;
    wire [3:0] lut_110_select = {
                             in_data[112],
                             in_data[56],
                             in_data[53],
                             in_data[72]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000000011110101;
    wire [3:0] lut_111_select = {
                             in_data[631],
                             in_data[707],
                             in_data[46],
                             in_data[118]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b0000000000101011;
    wire [3:0] lut_112_select = {
                             in_data[243],
                             in_data[216],
                             in_data[276],
                             in_data[206]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b1010101011111110;
    wire [3:0] lut_113_select = {
                             in_data[116],
                             in_data[449],
                             in_data[54],
                             in_data[103]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b0011001100100010;
    wire [3:0] lut_114_select = {
                             in_data[610],
                             in_data[14],
                             in_data[361],
                             in_data[274]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0011001100110011;
    wire [3:0] lut_115_select = {
                             in_data[763],
                             in_data[205],
                             in_data[267],
                             in_data[562]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b0100010001010101;
    wire [3:0] lut_116_select = {
                             in_data[548],
                             in_data[779],
                             in_data[531],
                             in_data[372]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b1011001110110011;
    wire [3:0] lut_117_select = {
                             in_data[670],
                             in_data[225],
                             in_data[634],
                             in_data[67]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1111111100100010;
    wire [3:0] lut_118_select = {
                             in_data[158],
                             in_data[756],
                             in_data[680],
                             in_data[78]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b0101010100000000;
    wire [3:0] lut_119_select = {
                             in_data[328],
                             in_data[421],
                             in_data[527],
                             in_data[90]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b0011000000110001;
    wire [3:0] lut_120_select = {
                             in_data[621],
                             in_data[309],
                             in_data[130],
                             in_data[701]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b0000000011111111;
    wire [3:0] lut_121_select = {
                             in_data[186],
                             in_data[460],
                             in_data[182],
                             in_data[607]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b0000100010101010;
    wire [3:0] lut_122_select = {
                             in_data[566],
                             in_data[48],
                             in_data[308],
                             in_data[241]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b1100111111001111;
    wire [3:0] lut_123_select = {
                             in_data[51],
                             in_data[272],
                             in_data[501],
                             in_data[474]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b1100110011001111;
    wire [3:0] lut_124_select = {
                             in_data[757],
                             in_data[188],
                             in_data[385],
                             in_data[52]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b0000111100000000;
    wire [3:0] lut_125_select = {
                             in_data[636],
                             in_data[535],
                             in_data[2],
                             in_data[195]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b1111111110100000;
    wire [3:0] lut_126_select = {
                             in_data[100],
                             in_data[244],
                             in_data[279],
                             in_data[326]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0001001100110011;
    wire [3:0] lut_127_select = {
                             in_data[177],
                             in_data[18],
                             in_data[355],
                             in_data[597]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b0101001001010101;
    wire [3:0] lut_128_select = {
                             in_data[271],
                             in_data[665],
                             in_data[128],
                             in_data[295]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b1111111111001110;
    wire [3:0] lut_129_select = {
                             in_data[741],
                             in_data[215],
                             in_data[626],
                             in_data[568]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b1101000011010000;
    wire [3:0] lut_130_select = {
                             in_data[57],
                             in_data[378],
                             in_data[704],
                             in_data[641]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b0101010101010101;
    wire [3:0] lut_131_select = {
                             in_data[364],
                             in_data[10],
                             in_data[31],
                             in_data[235]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b0101000101010001;
    wire [3:0] lut_132_select = {
                             in_data[644],
                             in_data[136],
                             in_data[466],
                             in_data[440]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0000000001011111;
    wire [3:0] lut_133_select = {
                             in_data[373],
                             in_data[110],
                             in_data[176],
                             in_data[482]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b1100111110001110;
    wire [3:0] lut_134_select = {
                             in_data[584],
                             in_data[685],
                             in_data[490],
                             in_data[723]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b0000000000010001;
    wire [3:0] lut_135_select = {
                             in_data[485],
                             in_data[559],
                             in_data[428],
                             in_data[102]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b0000111111111100;
    wire [3:0] lut_136_select = {
                             in_data[299],
                             in_data[119],
                             in_data[229],
                             in_data[503]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b0000000011110000;
    wire [3:0] lut_137_select = {
                             in_data[525],
                             in_data[327],
                             in_data[61],
                             in_data[60]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b0000000000000101;
    wire [3:0] lut_138_select = {
                             in_data[76],
                             in_data[511],
                             in_data[534],
                             in_data[75]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b0000000001000100;
    wire [3:0] lut_139_select = {
                             in_data[189],
                             in_data[506],
                             in_data[656],
                             in_data[137]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b0000000000010001;
    wire [3:0] lut_140_select = {
                             in_data[47],
                             in_data[16],
                             in_data[41],
                             in_data[497]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b0101010101000101;
    wire [3:0] lut_141_select = {
                             in_data[705],
                             in_data[601],
                             in_data[303],
                             in_data[443]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b1111000011111101;
    wire [3:0] lut_142_select = {
                             in_data[273],
                             in_data[38],
                             in_data[165],
                             in_data[765]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0000000000100010;
    wire [3:0] lut_143_select = {
                             in_data[611],
                             in_data[592],
                             in_data[304],
                             in_data[352]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b0000001000110011;
    wire [3:0] lut_144_select = {
                             in_data[157],
                             in_data[618],
                             in_data[403],
                             in_data[228]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1111111011111110;
    wire [3:0] lut_145_select = {
                             in_data[687],
                             in_data[745],
                             in_data[405],
                             in_data[771]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1010101010101010;
    wire [3:0] lut_146_select = {
                             in_data[781],
                             in_data[245],
                             in_data[234],
                             in_data[483]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0000000000000001;
    wire [3:0] lut_147_select = {
                             in_data[673],
                             in_data[367],
                             in_data[115],
                             in_data[742]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b0001001100000000;
    wire [3:0] lut_148_select = {
                             in_data[668],
                             in_data[747],
                             in_data[743],
                             in_data[365]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b1111101011111000;
    wire [3:0] lut_149_select = {
                             in_data[702],
                             in_data[353],
                             in_data[134],
                             in_data[174]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b0000000000010011;
    wire [3:0] lut_150_select = {
                             in_data[202],
                             in_data[36],
                             in_data[572],
                             in_data[604]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b0000000010101010;
    wire [3:0] lut_151_select = {
                             in_data[549],
                             in_data[389],
                             in_data[588],
                             in_data[407]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b0010001011101110;
    wire [3:0] lut_152_select = {
                             in_data[489],
                             in_data[576],
                             in_data[540],
                             in_data[297]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b0000000000010010;
    wire [3:0] lut_153_select = {
                             in_data[342],
                             in_data[602],
                             in_data[746],
                             in_data[713]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0001000000110000;
    wire [3:0] lut_154_select = {
                             in_data[193],
                             in_data[377],
                             in_data[415],
                             in_data[109]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b1010000010100001;
    wire [3:0] lut_155_select = {
                             in_data[418],
                             in_data[516],
                             in_data[366],
                             in_data[217]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b0010101010101110;
    wire [3:0] lut_156_select = {
                             in_data[620],
                             in_data[399],
                             in_data[435],
                             in_data[305]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b0000000000001110;
    wire [3:0] lut_157_select = {
                             in_data[508],
                             in_data[524],
                             in_data[334],
                             in_data[401]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b1000000011111101;
    wire [3:0] lut_158_select = {
                             in_data[467],
                             in_data[223],
                             in_data[80],
                             in_data[74]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b1111010111010101;
    wire [3:0] lut_159_select = {
                             in_data[33],
                             in_data[73],
                             in_data[363],
                             in_data[306]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b1111111111111011;
    wire [3:0] lut_160_select = {
                             in_data[512],
                             in_data[714],
                             in_data[347],
                             in_data[338]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b0000000001000100;
    wire [3:0] lut_161_select = {
                             in_data[429],
                             in_data[44],
                             in_data[151],
                             in_data[106]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1100000111000001;
    wire [3:0] lut_162_select = {
                             in_data[458],
                             in_data[567],
                             in_data[681],
                             in_data[310]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b1111001011110010;
    wire [3:0] lut_163_select = {
                             in_data[58],
                             in_data[722],
                             in_data[777],
                             in_data[740]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b1010101011111010;
    wire [3:0] lut_164_select = {
                             in_data[43],
                             in_data[716],
                             in_data[732],
                             in_data[266]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b0000111110101111;
    wire [3:0] lut_165_select = {
                             in_data[545],
                             in_data[184],
                             in_data[447],
                             in_data[316]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b1100110111001100;
    wire [3:0] lut_166_select = {
                             in_data[83],
                             in_data[412],
                             in_data[582],
                             in_data[63]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b1100101111001110;
    wire [3:0] lut_167_select = {
                             in_data[321],
                             in_data[499],
                             in_data[343],
                             in_data[275]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b0000000001010101;
    wire [3:0] lut_168_select = {
                             in_data[302],
                             in_data[42],
                             in_data[734],
                             in_data[689]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b1110110011111111;
    wire [3:0] lut_169_select = {
                             in_data[521],
                             in_data[675],
                             in_data[91],
                             in_data[614]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b0011000000110001;
    wire [3:0] lut_170_select = {
                             in_data[55],
                             in_data[8],
                             in_data[536],
                             in_data[758]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b1111111111111111;
    wire [3:0] lut_171_select = {
                             in_data[646],
                             in_data[281],
                             in_data[479],
                             in_data[669]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b0100010001001101;
    wire [3:0] lut_172_select = {
                             in_data[782],
                             in_data[718],
                             in_data[387],
                             in_data[652]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b1011000010110001;
    wire [3:0] lut_173_select = {
                             in_data[149],
                             in_data[290],
                             in_data[712],
                             in_data[551]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b0000000011011101;
    wire [3:0] lut_174_select = {
                             in_data[199],
                             in_data[392],
                             in_data[39],
                             in_data[214]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1111001111110011;
    wire [3:0] lut_175_select = {
                             in_data[82],
                             in_data[417],
                             in_data[348],
                             in_data[624]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b0000010100000001;
    wire [3:0] lut_176_select = {
                             in_data[724],
                             in_data[623],
                             in_data[236],
                             in_data[767]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b1110111011101110;
    wire [3:0] lut_177_select = {
                             in_data[169],
                             in_data[368],
                             in_data[737],
                             in_data[655]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b1111111110111010;
    wire [3:0] lut_178_select = {
                             in_data[411],
                             in_data[426],
                             in_data[21],
                             in_data[414]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b0101010111111111;
    wire [3:0] lut_179_select = {
                             in_data[237],
                             in_data[70],
                             in_data[84],
                             in_data[462]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b1111110011111111;
    wire [3:0] lut_180_select = {
                             in_data[181],
                             in_data[692],
                             in_data[543],
                             in_data[755]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b1001101100010001;
    wire [3:0] lut_181_select = {
                             in_data[207],
                             in_data[35],
                             in_data[380],
                             in_data[132]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b0000001100000011;
    wire [3:0] lut_182_select = {
                             in_data[251],
                             in_data[133],
                             in_data[156],
                             in_data[587]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b0000000000010001;
    wire [3:0] lut_183_select = {
                             in_data[654],
                             in_data[730],
                             in_data[627],
                             in_data[277]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b0011000101110101;
    wire [3:0] lut_184_select = {
                             in_data[768],
                             in_data[557],
                             in_data[264],
                             in_data[578]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b0000000000010001;
    wire [3:0] lut_185_select = {
                             in_data[79],
                             in_data[22],
                             in_data[619],
                             in_data[664]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b1010101010111010;
    wire [3:0] lut_186_select = {
                             in_data[81],
                             in_data[384],
                             in_data[3],
                             in_data[359]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b1100110011011111;
    wire [3:0] lut_187_select = {
                             in_data[632],
                             in_data[341],
                             in_data[484],
                             in_data[340]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b1010101110100010;
    wire [3:0] lut_188_select = {
                             in_data[456],
                             in_data[318],
                             in_data[198],
                             in_data[408]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b1011111111111010;
    wire [3:0] lut_189_select = {
                             in_data[187],
                             in_data[294],
                             in_data[731],
                             in_data[173]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b1111111111111010;
    wire [3:0] lut_190_select = {
                             in_data[269],
                             in_data[218],
                             in_data[441],
                             in_data[772]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b1111111010111010;
    wire [3:0] lut_191_select = {
                             in_data[329],
                             in_data[553],
                             in_data[555],
                             in_data[349]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b0101110001001100;
    wire [3:0] lut_192_select = {
                             in_data[672],
                             in_data[469],
                             in_data[433],
                             in_data[579]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b1111001011110011;
    wire [3:0] lut_193_select = {
                             in_data[252],
                             in_data[312],
                             in_data[221],
                             in_data[25]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0100110000001111;
    wire [3:0] lut_194_select = {
                             in_data[268],
                             in_data[344],
                             in_data[98],
                             in_data[505]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b0001110100001100;
    wire [3:0] lut_195_select = {
                             in_data[542],
                             in_data[370],
                             in_data[526],
                             in_data[651]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b1111101111110000;
    wire [3:0] lut_196_select = {
                             in_data[528],
                             in_data[488],
                             in_data[285],
                             in_data[460]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b1111111100001100;
    wire [3:0] lut_197_select = {
                             in_data[539],
                             in_data[649],
                             in_data[179],
                             in_data[224]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b1001100110011001;
    wire [3:0] lut_198_select = {
                             in_data[374],
                             in_data[30],
                             in_data[541],
                             in_data[538]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b0000001100000011;
    wire [3:0] lut_199_select = {
                             in_data[643],
                             in_data[208],
                             in_data[298],
                             in_data[0]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b0000001000000011;
    wire [3:0] lut_200_select = {
                             in_data[737],
                             in_data[370],
                             in_data[709],
                             in_data[307]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b0000000100000001;
    wire [3:0] lut_201_select = {
                             in_data[588],
                             in_data[395],
                             in_data[444],
                             in_data[500]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b0000001000110011;
    wire [3:0] lut_202_select = {
                             in_data[496],
                             in_data[343],
                             in_data[442],
                             in_data[481]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b0000000011000011;
    wire [3:0] lut_203_select = {
                             in_data[581],
                             in_data[691],
                             in_data[398],
                             in_data[14]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b0000110000001111;
    wire [3:0] lut_204_select = {
                             in_data[663],
                             in_data[459],
                             in_data[302],
                             in_data[59]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b1111111111111100;
    wire [3:0] lut_205_select = {
                             in_data[260],
                             in_data[345],
                             in_data[733],
                             in_data[363]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b1100110011101110;
    wire [3:0] lut_206_select = {
                             in_data[308],
                             in_data[2],
                             in_data[620],
                             in_data[704]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b1111110111111100;
    wire [3:0] lut_207_select = {
                             in_data[251],
                             in_data[68],
                             in_data[542],
                             in_data[665]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1111111111111110;
    wire [3:0] lut_208_select = {
                             in_data[611],
                             in_data[124],
                             in_data[299],
                             in_data[283]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b0101111101011111;
    wire [3:0] lut_209_select = {
                             in_data[755],
                             in_data[408],
                             in_data[169],
                             in_data[599]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b0000000011111111;
    wire [3:0] lut_210_select = {
                             in_data[400],
                             in_data[672],
                             in_data[636],
                             in_data[449]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b0000000011001111;
    wire [3:0] lut_211_select = {
                             in_data[323],
                             in_data[674],
                             in_data[607],
                             in_data[61]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b0000111000001110;
    wire [3:0] lut_212_select = {
                             in_data[7],
                             in_data[262],
                             in_data[623],
                             in_data[465]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b1110010001000100;
    wire [3:0] lut_213_select = {
                             in_data[632],
                             in_data[202],
                             in_data[324],
                             in_data[580]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1111111111111110;
    wire [3:0] lut_214_select = {
                             in_data[751],
                             in_data[432],
                             in_data[446],
                             in_data[77]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b1101110011111100;
    wire [3:0] lut_215_select = {
                             in_data[411],
                             in_data[319],
                             in_data[692],
                             in_data[243]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b0100010011100111;
    wire [3:0] lut_216_select = {
                             in_data[234],
                             in_data[472],
                             in_data[693],
                             in_data[575]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b1111111111101110;
    wire [3:0] lut_217_select = {
                             in_data[624],
                             in_data[420],
                             in_data[687],
                             in_data[390]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b0000001100000011;
    wire [3:0] lut_218_select = {
                             in_data[140],
                             in_data[711],
                             in_data[768],
                             in_data[605]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b1100111111001101;
    wire [3:0] lut_219_select = {
                             in_data[8],
                             in_data[186],
                             in_data[342],
                             in_data[326]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b0000000100000001;
    wire [3:0] lut_220_select = {
                             in_data[166],
                             in_data[119],
                             in_data[382],
                             in_data[551]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b1010101011111010;
    wire [3:0] lut_221_select = {
                             in_data[195],
                             in_data[419],
                             in_data[476],
                             in_data[367]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b0011001100110011;
    wire [3:0] lut_222_select = {
                             in_data[82],
                             in_data[144],
                             in_data[397],
                             in_data[200]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1111111111111010;
    wire [3:0] lut_223_select = {
                             in_data[192],
                             in_data[719],
                             in_data[180],
                             in_data[402]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b0001010101010101;
    wire [3:0] lut_224_select = {
                             in_data[702],
                             in_data[724],
                             in_data[600],
                             in_data[656]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b0000111100001111;
    wire [3:0] lut_225_select = {
                             in_data[546],
                             in_data[601],
                             in_data[467],
                             in_data[477]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1011101110111011;
    wire [3:0] lut_226_select = {
                             in_data[583],
                             in_data[586],
                             in_data[682],
                             in_data[536]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b1110111011101110;
    wire [3:0] lut_227_select = {
                             in_data[593],
                             in_data[645],
                             in_data[214],
                             in_data[358]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b0001001100010011;
    wire [3:0] lut_228_select = {
                             in_data[749],
                             in_data[130],
                             in_data[659],
                             in_data[286]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b0000000000110000;
    wire [3:0] lut_229_select = {
                             in_data[315],
                             in_data[653],
                             in_data[641],
                             in_data[313]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b1111111111101111;
    wire [3:0] lut_230_select = {
                             in_data[132],
                             in_data[207],
                             in_data[483],
                             in_data[94]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b0111001111110011;
    wire [3:0] lut_231_select = {
                             in_data[280],
                             in_data[594],
                             in_data[517],
                             in_data[695]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b0001000100010001;
    wire [3:0] lut_232_select = {
                             in_data[560],
                             in_data[87],
                             in_data[531],
                             in_data[573]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b1111000001000100;
    wire [3:0] lut_233_select = {
                             in_data[353],
                             in_data[184],
                             in_data[708],
                             in_data[41]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b1111101111111011;
    wire [3:0] lut_234_select = {
                             in_data[730],
                             in_data[613],
                             in_data[438],
                             in_data[90]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b1010101010101010;
    wire [3:0] lut_235_select = {
                             in_data[756],
                             in_data[175],
                             in_data[121],
                             in_data[384]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b0101000001010101;
    wire [3:0] lut_236_select = {
                             in_data[242],
                             in_data[230],
                             in_data[713],
                             in_data[310]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b0101010100000101;
    wire [3:0] lut_237_select = {
                             in_data[222],
                             in_data[379],
                             in_data[752],
                             in_data[559]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b1111111110101010;
    wire [3:0] lut_238_select = {
                             in_data[712],
                             in_data[80],
                             in_data[759],
                             in_data[328]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0000000001010101;
    wire [3:0] lut_239_select = {
                             in_data[248],
                             in_data[23],
                             in_data[783],
                             in_data[375]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b1011111110101010;
    wire [3:0] lut_240_select = {
                             in_data[114],
                             in_data[503],
                             in_data[673],
                             in_data[229]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b1111111111001000;
    wire [3:0] lut_241_select = {
                             in_data[489],
                             in_data[361],
                             in_data[431],
                             in_data[316]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b1010111110101111;
    wire [3:0] lut_242_select = {
                             in_data[777],
                             in_data[552],
                             in_data[4],
                             in_data[368]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b1010101011101010;
    wire [3:0] lut_243_select = {
                             in_data[64],
                             in_data[291],
                             in_data[85],
                             in_data[596]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b0000010001000101;
    wire [3:0] lut_244_select = {
                             in_data[18],
                             in_data[137],
                             in_data[340],
                             in_data[78]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b1111111011101110;
    wire [3:0] lut_245_select = {
                             in_data[521],
                             in_data[527],
                             in_data[176],
                             in_data[354]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b1110111111101111;
    wire [3:0] lut_246_select = {
                             in_data[167],
                             in_data[603],
                             in_data[341],
                             in_data[344]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b0000000000000001;
    wire [3:0] lut_247_select = {
                             in_data[360],
                             in_data[231],
                             in_data[331],
                             in_data[272]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b0001000100010001;
    wire [3:0] lut_248_select = {
                             in_data[757],
                             in_data[51],
                             in_data[661],
                             in_data[161]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b0000010000001111;
    wire [3:0] lut_249_select = {
                             in_data[462],
                             in_data[428],
                             in_data[233],
                             in_data[98]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b1111001111110011;
    wire [3:0] lut_250_select = {
                             in_data[281],
                             in_data[136],
                             in_data[203],
                             in_data[226]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b1110111011101110;
    wire [3:0] lut_251_select = {
                             in_data[615],
                             in_data[639],
                             in_data[97],
                             in_data[131]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b1011001100000000;
    wire [3:0] lut_252_select = {
                             in_data[433],
                             in_data[574],
                             in_data[235],
                             in_data[764]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b1110110011101100;
    wire [3:0] lut_253_select = {
                             in_data[11],
                             in_data[122],
                             in_data[681],
                             in_data[213]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b0000000011111110;
    wire [3:0] lut_254_select = {
                             in_data[710],
                             in_data[545],
                             in_data[587],
                             in_data[105]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b0010101000101010;
    wire [3:0] lut_255_select = {
                             in_data[1],
                             in_data[279],
                             in_data[170],
                             in_data[471]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b0000000000010000;
    wire [3:0] lut_256_select = {
                             in_data[732],
                             in_data[540],
                             in_data[745],
                             in_data[422]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b1111111111111100;
    wire [3:0] lut_257_select = {
                             in_data[417],
                             in_data[501],
                             in_data[727],
                             in_data[701]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b0010000001011111;
    wire [3:0] lut_258_select = {
                             in_data[598],
                             in_data[256],
                             in_data[690],
                             in_data[434]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b0000000000000011;
    wire [3:0] lut_259_select = {
                             in_data[102],
                             in_data[565],
                             in_data[160],
                             in_data[21]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b1111101011111010;
    wire [3:0] lut_260_select = {
                             in_data[115],
                             in_data[482],
                             in_data[533],
                             in_data[470]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b1011001111110011;
    wire [3:0] lut_261_select = {
                             in_data[734],
                             in_data[748],
                             in_data[406],
                             in_data[52]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b0010000011110011;
    wire [3:0] lut_262_select = {
                             in_data[775],
                             in_data[590],
                             in_data[289],
                             in_data[418]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b0000101100001010;
    wire [3:0] lut_263_select = {
                             in_data[750],
                             in_data[512],
                             in_data[414],
                             in_data[321]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b0101111101011111;
    wire [3:0] lut_264_select = {
                             in_data[47],
                             in_data[264],
                             in_data[771],
                             in_data[346]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b0000000001010000;
    wire [3:0] lut_265_select = {
                             in_data[766],
                             in_data[487],
                             in_data[731],
                             in_data[221]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1110110011111100;
    wire [3:0] lut_266_select = {
                             in_data[95],
                             in_data[325],
                             in_data[255],
                             in_data[365]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b0000000011111111;
    wire [3:0] lut_267_select = {
                             in_data[513],
                             in_data[421],
                             in_data[60],
                             in_data[424]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1000000011111101;
    wire [3:0] lut_268_select = {
                             in_data[339],
                             in_data[445],
                             in_data[104],
                             in_data[381]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0100010100000100;
    wire [3:0] lut_269_select = {
                             in_data[296],
                             in_data[668],
                             in_data[74],
                             in_data[582]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b1111111111001110;
    wire [3:0] lut_270_select = {
                             in_data[125],
                             in_data[627],
                             in_data[413],
                             in_data[201]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b1111111110101010;
    wire [3:0] lut_271_select = {
                             in_data[507],
                             in_data[168],
                             in_data[88],
                             in_data[436]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b0011010011111110;
    wire [3:0] lut_272_select = {
                             in_data[362],
                             in_data[484],
                             in_data[485],
                             in_data[287]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b0000111100001101;
    wire [3:0] lut_273_select = {
                             in_data[84],
                             in_data[120],
                             in_data[86],
                             in_data[683]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b0000110000001110;
    wire [3:0] lut_274_select = {
                             in_data[633],
                             in_data[333],
                             in_data[427],
                             in_data[781]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b0000010100000101;
    wire [3:0] lut_275_select = {
                             in_data[334],
                             in_data[250],
                             in_data[3],
                             in_data[405]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b1010111011101110;
    wire [3:0] lut_276_select = {
                             in_data[336],
                             in_data[73],
                             in_data[178],
                             in_data[621]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b0000000000110011;
    wire [3:0] lut_277_select = {
                             in_data[212],
                             in_data[20],
                             in_data[312],
                             in_data[29]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b0101010101010101;
    wire [3:0] lut_278_select = {
                             in_data[616],
                             in_data[698],
                             in_data[650],
                             in_data[371]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b0000101100000011;
    wire [3:0] lut_279_select = {
                             in_data[50],
                             in_data[274],
                             in_data[416],
                             in_data[776]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b0001000000110000;
    wire [3:0] lut_280_select = {
                             in_data[778],
                             in_data[456],
                             in_data[172],
                             in_data[564]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b1111111111111100;
    wire [3:0] lut_281_select = {
                             in_data[505],
                             in_data[123],
                             in_data[780],
                             in_data[25]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b0001000011110001;
    wire [3:0] lut_282_select = {
                             in_data[563],
                             in_data[739],
                             in_data[211],
                             in_data[118]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b0000101000001111;
    wire [3:0] lut_283_select = {
                             in_data[450],
                             in_data[352],
                             in_data[34],
                             in_data[349]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b1011001100000001;
    wire [3:0] lut_284_select = {
                             in_data[440],
                             in_data[523],
                             in_data[566],
                             in_data[666]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b1111111111110001;
    wire [3:0] lut_285_select = {
                             in_data[686],
                             in_data[164],
                             in_data[141],
                             in_data[265]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b0000000011111011;
    wire [3:0] lut_286_select = {
                             in_data[454],
                             in_data[145],
                             in_data[139],
                             in_data[729]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b0011000011110100;
    wire [3:0] lut_287_select = {
                             in_data[425],
                             in_data[156],
                             in_data[181],
                             in_data[58]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b0001010100010001;
    wire [3:0] lut_288_select = {
                             in_data[5],
                             in_data[117],
                             in_data[153],
                             in_data[572]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b0101010101010001;
    wire [3:0] lut_289_select = {
                             in_data[27],
                             in_data[753],
                             in_data[19],
                             in_data[721]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b1000101011101110;
    wire [3:0] lut_290_select = {
                             in_data[72],
                             in_data[17],
                             in_data[628],
                             in_data[736]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b0000010100000101;
    wire [3:0] lut_291_select = {
                             in_data[171],
                             in_data[608],
                             in_data[716],
                             in_data[275]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b0000000000000100;
    wire [3:0] lut_292_select = {
                             in_data[79],
                             in_data[747],
                             in_data[56],
                             in_data[311]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b0101010001010100;
    wire [3:0] lut_293_select = {
                             in_data[22],
                             in_data[399],
                             in_data[671],
                             in_data[725]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1111111100001100;
    wire [3:0] lut_294_select = {
                             in_data[189],
                             in_data[148],
                             in_data[187],
                             in_data[16]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b0100010011111111;
    wire [3:0] lut_295_select = {
                             in_data[490],
                             in_data[675],
                             in_data[65],
                             in_data[609]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b1111110100100000;
    wire [3:0] lut_296_select = {
                             in_data[544],
                             in_data[706],
                             in_data[654],
                             in_data[271]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b1111111100001110;
    wire [3:0] lut_297_select = {
                             in_data[149],
                             in_data[389],
                             in_data[614],
                             in_data[494]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b1111110111011101;
    wire [3:0] lut_298_select = {
                             in_data[236],
                             in_data[534],
                             in_data[304],
                             in_data[543]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b1111111110111010;
    wire [3:0] lut_299_select = {
                             in_data[205],
                             in_data[670],
                             in_data[107],
                             in_data[769]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b0000000100000001;
    wire [3:0] lut_300_select = {
                             in_data[642],
                             in_data[746],
                             in_data[741],
                             in_data[129]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b0010001100000010;
    wire [3:0] lut_301_select = {
                             in_data[480],
                             in_data[526],
                             in_data[76],
                             in_data[410]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b0000010001001101;
    wire [3:0] lut_302_select = {
                             in_data[297],
                             in_data[451],
                             in_data[570],
                             in_data[423]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b1010101110101011;
    wire [3:0] lut_303_select = {
                             in_data[644],
                             in_data[634],
                             in_data[348],
                             in_data[282]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b0000000000001100;
    wire [3:0] lut_304_select = {
                             in_data[71],
                             in_data[415],
                             in_data[232],
                             in_data[75]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b0000000000000011;
    wire [3:0] lut_305_select = {
                             in_data[502],
                             in_data[396],
                             in_data[219],
                             in_data[32]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b1010101110101011;
    wire [3:0] lut_306_select = {
                             in_data[48],
                             in_data[401],
                             in_data[474],
                             in_data[152]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b1111000010101011;
    wire [3:0] lut_307_select = {
                             in_data[514],
                             in_data[508],
                             in_data[782],
                             in_data[293]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b0000000000000011;
    wire [3:0] lut_308_select = {
                             in_data[330],
                             in_data[103],
                             in_data[254],
                             in_data[33]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b0001000000010000;
    wire [3:0] lut_309_select = {
                             in_data[618],
                             in_data[237],
                             in_data[159],
                             in_data[347]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b1111111111110110;
    wire [3:0] lut_310_select = {
                             in_data[217],
                             in_data[604],
                             in_data[651],
                             in_data[567]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b1010101010101010;
    wire [3:0] lut_311_select = {
                             in_data[754],
                             in_data[10],
                             in_data[700],
                             in_data[655]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1010000010101110;
    wire [3:0] lut_312_select = {
                             in_data[322],
                             in_data[715],
                             in_data[364],
                             in_data[327]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b1111111100000100;
    wire [3:0] lut_313_select = {
                             in_data[412],
                             in_data[667],
                             in_data[252],
                             in_data[393]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b0000000011101110;
    wire [3:0] lut_314_select = {
                             in_data[185],
                             in_data[763],
                             in_data[292],
                             in_data[295]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b1111011111110100;
    wire [3:0] lut_315_select = {
                             in_data[288],
                             in_data[177],
                             in_data[155],
                             in_data[106]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b1000101010000011;
    wire [3:0] lut_316_select = {
                             in_data[597],
                             in_data[509],
                             in_data[458],
                             in_data[557]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b0000000000100011;
    wire [3:0] lut_317_select = {
                             in_data[558],
                             in_data[699],
                             in_data[678],
                             in_data[15]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0000010100000000;
    wire [3:0] lut_318_select = {
                             in_data[548],
                             in_data[705],
                             in_data[617],
                             in_data[738]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b1100110000000011;
    wire [3:0] lut_319_select = {
                             in_data[244],
                             in_data[491],
                             in_data[463],
                             in_data[391]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b0101000101010101;
    wire [3:0] lut_320_select = {
                             in_data[329],
                             in_data[740],
                             in_data[525],
                             in_data[162]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0000000001010101;
    wire [3:0] lut_321_select = {
                             in_data[383],
                             in_data[225],
                             in_data[475],
                             in_data[270]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b1100110011001100;
    wire [3:0] lut_322_select = {
                             in_data[720],
                             in_data[301],
                             in_data[294],
                             in_data[108]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b1111110011001100;
    wire [3:0] lut_323_select = {
                             in_data[261],
                             in_data[183],
                             in_data[239],
                             in_data[519]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b0100010001010101;
    wire [3:0] lut_324_select = {
                             in_data[437],
                             in_data[647],
                             in_data[591],
                             in_data[714]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b1111111100000000;
    wire [3:0] lut_325_select = {
                             in_data[569],
                             in_data[257],
                             in_data[116],
                             in_data[758]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b0000000010110010;
    wire [3:0] lut_326_select = {
                             in_data[664],
                             in_data[498],
                             in_data[703],
                             in_data[13]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b1010101010101110;
    wire [3:0] lut_327_select = {
                             in_data[635],
                             in_data[637],
                             in_data[529],
                             in_data[157]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b1111111111110000;
    wire [3:0] lut_328_select = {
                             in_data[499],
                             in_data[246],
                             in_data[45],
                             in_data[774]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b0000101000001111;
    wire [3:0] lut_329_select = {
                             in_data[435],
                             in_data[228],
                             in_data[113],
                             in_data[259]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b1111111101000101;
    wire [3:0] lut_330_select = {
                             in_data[300],
                             in_data[109],
                             in_data[28],
                             in_data[602]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b0000000000000101;
    wire [3:0] lut_331_select = {
                             in_data[535],
                             in_data[133],
                             in_data[83],
                             in_data[154]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b0101101011111010;
    wire [3:0] lut_332_select = {
                             in_data[696],
                             in_data[457],
                             in_data[760],
                             in_data[515]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b1111110111111110;
    wire [3:0] lut_333_select = {
                             in_data[314],
                             in_data[267],
                             in_data[742],
                             in_data[332]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b0000000000001100;
    wire [3:0] lut_334_select = {
                             in_data[443],
                             in_data[592],
                             in_data[268],
                             in_data[42]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0011001100110011;
    wire [3:0] lut_335_select = {
                             in_data[357],
                             in_data[44],
                             in_data[158],
                             in_data[657]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b0000010100000101;
    wire [3:0] lut_336_select = {
                             in_data[726],
                             in_data[464],
                             in_data[55],
                             in_data[638]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b1110111111101110;
    wire [3:0] lut_337_select = {
                             in_data[67],
                             in_data[240],
                             in_data[218],
                             in_data[306]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b1100110011001101;
    wire [3:0] lut_338_select = {
                             in_data[35],
                             in_data[595],
                             in_data[473],
                             in_data[335]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b0101010111001111;
    wire [3:0] lut_339_select = {
                             in_data[430],
                             in_data[767],
                             in_data[81],
                             in_data[182]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b0111100001010000;
    wire [3:0] lut_340_select = {
                             in_data[143],
                             in_data[626],
                             in_data[93],
                             in_data[355]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b1111101011111111;
    wire [3:0] lut_341_select = {
                             in_data[761],
                             in_data[676],
                             in_data[337],
                             in_data[735]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b0000000000110011;
    wire [3:0] lut_342_select = {
                             in_data[684],
                             in_data[111],
                             in_data[165],
                             in_data[258]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b0010001000100110;
    wire [3:0] lut_343_select = {
                             in_data[138],
                             in_data[223],
                             in_data[466],
                             in_data[351]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1111101011110010;
    wire [3:0] lut_344_select = {
                             in_data[173],
                             in_data[492],
                             in_data[190],
                             in_data[100]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b0000000000100011;
    wire [3:0] lut_345_select = {
                             in_data[338],
                             in_data[447],
                             in_data[269],
                             in_data[669]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b0000001100000011;
    wire [3:0] lut_346_select = {
                             in_data[779],
                             in_data[478],
                             in_data[403],
                             in_data[53]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b0001000100000001;
    wire [3:0] lut_347_select = {
                             in_data[532],
                             in_data[550],
                             in_data[562],
                             in_data[495]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0000000000000001;
    wire [3:0] lut_348_select = {
                             in_data[772],
                             in_data[537],
                             in_data[247],
                             in_data[204]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b0000001100000011;
    wire [3:0] lut_349_select = {
                             in_data[448],
                             in_data[273],
                             in_data[522],
                             in_data[62]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b0000000000000000;
    wire [3:0] lut_350_select = {
                             in_data[197],
                             in_data[479],
                             in_data[194],
                             in_data[63]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b1100111101001100;
    wire [3:0] lut_351_select = {
                             in_data[629],
                             in_data[640],
                             in_data[193],
                             in_data[622]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b0000000011010101;
    wire [3:0] lut_352_select = {
                             in_data[554],
                             in_data[762],
                             in_data[163],
                             in_data[43]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b0011000000110000;
    wire [3:0] lut_353_select = {
                             in_data[658],
                             in_data[290],
                             in_data[278],
                             in_data[728]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b0000000000000011;
    wire [3:0] lut_354_select = {
                             in_data[146],
                             in_data[571],
                             in_data[96],
                             in_data[773]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b0001000001010000;
    wire [3:0] lut_355_select = {
                             in_data[579],
                             in_data[409],
                             in_data[46],
                             in_data[612]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b1101010111010101;
    wire [3:0] lut_356_select = {
                             in_data[134],
                             in_data[40],
                             in_data[126],
                             in_data[493]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b0000010100000000;
    wire [3:0] lut_357_select = {
                             in_data[429],
                             in_data[99],
                             in_data[198],
                             in_data[277]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b0000110111001100;
    wire [3:0] lut_358_select = {
                             in_data[376],
                             in_data[707],
                             in_data[606],
                             in_data[516]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b1111111101010000;
    wire [3:0] lut_359_select = {
                             in_data[439],
                             in_data[388],
                             in_data[392],
                             in_data[518]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b1111101011111100;
    wire [3:0] lut_360_select = {
                             in_data[630],
                             in_data[151],
                             in_data[373],
                             in_data[589]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b1110110011101110;
    wire [3:0] lut_361_select = {
                             in_data[245],
                             in_data[577],
                             in_data[576],
                             in_data[66]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b0010011101010000;
    wire [3:0] lut_362_select = {
                             in_data[378],
                             in_data[206],
                             in_data[49],
                             in_data[404]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b0101000011010101;
    wire [3:0] lut_363_select = {
                             in_data[372],
                             in_data[524],
                             in_data[646],
                             in_data[276]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b0101000001010101;
    wire [3:0] lut_364_select = {
                             in_data[350],
                             in_data[619],
                             in_data[238],
                             in_data[677]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b1100111100001100;
    wire [3:0] lut_365_select = {
                             in_data[506],
                             in_data[369],
                             in_data[553],
                             in_data[12]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b0000000000000001;
    wire [3:0] lut_366_select = {
                             in_data[662],
                             in_data[568],
                             in_data[511],
                             in_data[150]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b1111111101010101;
    wire [3:0] lut_367_select = {
                             in_data[744],
                             in_data[284],
                             in_data[585],
                             in_data[549]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b1111110011111100;
    wire [3:0] lut_368_select = {
                             in_data[452],
                             in_data[679],
                             in_data[356],
                             in_data[561]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b1111111111111100;
    wire [3:0] lut_369_select = {
                             in_data[317],
                             in_data[770],
                             in_data[303],
                             in_data[722]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b1111111111101110;
    wire [3:0] lut_370_select = {
                             in_data[625],
                             in_data[216],
                             in_data[101],
                             in_data[743]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b1111111111101110;
    wire [3:0] lut_371_select = {
                             in_data[263],
                             in_data[685],
                             in_data[249],
                             in_data[220]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b0001000101010101;
    wire [3:0] lut_372_select = {
                             in_data[128],
                             in_data[504],
                             in_data[556],
                             in_data[127]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b0000000001000100;
    wire [3:0] lut_373_select = {
                             in_data[469],
                             in_data[57],
                             in_data[241],
                             in_data[578]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b0101111100000000;
    wire [3:0] lut_374_select = {
                             in_data[209],
                             in_data[110],
                             in_data[253],
                             in_data[631]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b1111111111111010;
    wire [3:0] lut_375_select = {
                             in_data[407],
                             in_data[689],
                             in_data[199],
                             in_data[359]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b0011001011110011;
    wire [3:0] lut_376_select = {
                             in_data[135],
                             in_data[530],
                             in_data[320],
                             in_data[652]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b1111111111110011;
    wire [3:0] lut_377_select = {
                             in_data[70],
                             in_data[305],
                             in_data[486],
                             in_data[36]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b1111111111111111;
    wire [3:0] lut_378_select = {
                             in_data[309],
                             in_data[227],
                             in_data[39],
                             in_data[394]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1111111101010101;
    wire [3:0] lut_379_select = {
                             in_data[92],
                             in_data[112],
                             in_data[26],
                             in_data[453]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b1111000011110111;
    wire [3:0] lut_380_select = {
                             in_data[497],
                             in_data[717],
                             in_data[468],
                             in_data[366]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b0000000010101010;
    wire [3:0] lut_381_select = {
                             in_data[387],
                             in_data[69],
                             in_data[6],
                             in_data[266]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b0110111101001111;
    wire [3:0] lut_382_select = {
                             in_data[91],
                             in_data[210],
                             in_data[441],
                             in_data[174]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b0101000101010001;
    wire [3:0] lut_383_select = {
                             in_data[24],
                             in_data[680],
                             in_data[191],
                             in_data[215]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0000001100000011;
    wire [3:0] lut_384_select = {
                             in_data[54],
                             in_data[385],
                             in_data[694],
                             in_data[31]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b0011001100000000;
    wire [3:0] lut_385_select = {
                             in_data[461],
                             in_data[520],
                             in_data[555],
                             in_data[547]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b0000000011001100;
    wire [3:0] lut_386_select = {
                             in_data[723],
                             in_data[142],
                             in_data[510],
                             in_data[648]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b0111000011110010;
    wire [3:0] lut_387_select = {
                             in_data[765],
                             in_data[455],
                             in_data[386],
                             in_data[147]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b1100110011001100;
    wire [3:0] lut_388_select = {
                             in_data[9],
                             in_data[196],
                             in_data[380],
                             in_data[318]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b1100000011000001;
    wire [3:0] lut_389_select = {
                             in_data[584],
                             in_data[688],
                             in_data[610],
                             in_data[426]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b1111111111111110;
    wire [3:0] lut_390_select = {
                             in_data[697],
                             in_data[38],
                             in_data[89],
                             in_data[37]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b0100010101011101;
    wire [3:0] lut_391_select = {
                             in_data[188],
                             in_data[660],
                             in_data[718],
                             in_data[377]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b1111111101010100;
    wire [3:0] lut_392_select = {
                             in_data[124],
                             in_data[442],
                             in_data[771],
                             in_data[305]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b1111101011111010;
    wire [3:0] lut_393_select = {
                             in_data[9],
                             in_data[681],
                             in_data[212],
                             in_data[685]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b0001001100110001;
    wire [3:0] lut_394_select = {
                             in_data[203],
                             in_data[302],
                             in_data[317],
                             in_data[652]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b1111111100000000;
    wire [3:0] lut_395_select = {
                             in_data[570],
                             in_data[206],
                             in_data[701],
                             in_data[179]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b0000000011111100;
    wire [3:0] lut_396_select = {
                             in_data[370],
                             in_data[304],
                             in_data[323],
                             in_data[25]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b1010101010101010;
    wire [3:0] lut_397_select = {
                             in_data[475],
                             in_data[684],
                             in_data[243],
                             in_data[293]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b1111111111111100;
    wire [3:0] lut_398_select = {
                             in_data[444],
                             in_data[457],
                             in_data[396],
                             in_data[64]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b1010111100100010;
    wire [3:0] lut_399_select = {
                             in_data[375],
                             in_data[640],
                             in_data[176],
                             in_data[249]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b0010001010101010;
    wire [3:0] lut_400_select = {
                             in_data[752],
                             in_data[578],
                             in_data[708],
                             in_data[428]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b0001010100000001;
    wire [3:0] lut_401_select = {
                             in_data[218],
                             in_data[178],
                             in_data[310],
                             in_data[592]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b0000000100000000;
    wire [3:0] lut_402_select = {
                             in_data[463],
                             in_data[72],
                             in_data[92],
                             in_data[193]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b0011001100110011;
    wire [3:0] lut_403_select = {
                             in_data[11],
                             in_data[773],
                             in_data[403],
                             in_data[362]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b1010111110001111;
    wire [3:0] lut_404_select = {
                             in_data[774],
                             in_data[658],
                             in_data[433],
                             in_data[474]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b0000000011011101;
    wire [3:0] lut_405_select = {
                             in_data[192],
                             in_data[778],
                             in_data[605],
                             in_data[348]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0101010101010101;
    wire [3:0] lut_406_select = {
                             in_data[665],
                             in_data[779],
                             in_data[476],
                             in_data[453]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b0101110100000101;
    wire [3:0] lut_407_select = {
                             in_data[219],
                             in_data[99],
                             in_data[223],
                             in_data[430]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b0000001100000011;
    wire [3:0] lut_408_select = {
                             in_data[32],
                             in_data[568],
                             in_data[422],
                             in_data[730]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b0000010100001111;
    wire [3:0] lut_409_select = {
                             in_data[682],
                             in_data[445],
                             in_data[59],
                             in_data[407]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b0000000100000001;
    wire [3:0] lut_410_select = {
                             in_data[381],
                             in_data[165],
                             in_data[397],
                             in_data[316]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b0010001110101010;
    wire [3:0] lut_411_select = {
                             in_data[341],
                             in_data[123],
                             in_data[542],
                             in_data[290]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b0101010100000100;
    wire [3:0] lut_412_select = {
                             in_data[324],
                             in_data[735],
                             in_data[523],
                             in_data[569]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b1010101011111111;
    wire [3:0] lut_413_select = {
                             in_data[291],
                             in_data[10],
                             in_data[47],
                             in_data[455]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0000001100000011;
    wire [3:0] lut_414_select = {
                             in_data[352],
                             in_data[609],
                             in_data[152],
                             in_data[745]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b0001010100000000;
    wire [3:0] lut_415_select = {
                             in_data[320],
                             in_data[454],
                             in_data[432],
                             in_data[535]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b0101010100000000;
    wire [3:0] lut_416_select = {
                             in_data[657],
                             in_data[17],
                             in_data[618],
                             in_data[285]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b1111111100000100;
    wire [3:0] lut_417_select = {
                             in_data[413],
                             in_data[649],
                             in_data[71],
                             in_data[734]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b0011001100010001;
    wire [3:0] lut_418_select = {
                             in_data[502],
                             in_data[252],
                             in_data[549],
                             in_data[547]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b0000110000001111;
    wire [3:0] lut_419_select = {
                             in_data[180],
                             in_data[580],
                             in_data[334],
                             in_data[195]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b0001000001010000;
    wire [3:0] lut_420_select = {
                             in_data[229],
                             in_data[402],
                             in_data[629],
                             in_data[473]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b0000000001010101;
    wire [3:0] lut_421_select = {
                             in_data[183],
                             in_data[142],
                             in_data[31],
                             in_data[283]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b0010101000101010;
    wire [3:0] lut_422_select = {
                             in_data[8],
                             in_data[115],
                             in_data[146],
                             in_data[354]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b1101110111001101;
    wire [3:0] lut_423_select = {
                             in_data[417],
                             in_data[230],
                             in_data[276],
                             in_data[372]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b0000000000010001;
    wire [3:0] lut_424_select = {
                             in_data[594],
                             in_data[644],
                             in_data[664],
                             in_data[621]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b1101010111110101;
    wire [3:0] lut_425_select = {
                             in_data[571],
                             in_data[356],
                             in_data[676],
                             in_data[349]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b1111111110111011;
    wire [3:0] lut_426_select = {
                             in_data[257],
                             in_data[106],
                             in_data[458],
                             in_data[744]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b0101010111010101;
    wire [3:0] lut_427_select = {
                             in_data[438],
                             in_data[704],
                             in_data[662],
                             in_data[427]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b1111111111111100;
    wire [3:0] lut_428_select = {
                             in_data[687],
                             in_data[632],
                             in_data[250],
                             in_data[698]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b0000010001001100;
    wire [3:0] lut_429_select = {
                             in_data[494],
                             in_data[525],
                             in_data[627],
                             in_data[171]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b0011001000110011;
    wire [3:0] lut_430_select = {
                             in_data[521],
                             in_data[137],
                             in_data[418],
                             in_data[747]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b1111010111110000;
    wire [3:0] lut_431_select = {
                             in_data[429],
                             in_data[610],
                             in_data[782],
                             in_data[220]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b0000100010001110;
    wire [3:0] lut_432_select = {
                             in_data[742],
                             in_data[529],
                             in_data[272],
                             in_data[69]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b0101010101010101;
    wire [3:0] lut_433_select = {
                             in_data[566],
                             in_data[364],
                             in_data[18],
                             in_data[481]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b0000111100001111;
    wire [3:0] lut_434_select = {
                             in_data[661],
                             in_data[490],
                             in_data[154],
                             in_data[638]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b0000111100001100;
    wire [3:0] lut_435_select = {
                             in_data[14],
                             in_data[695],
                             in_data[189],
                             in_data[26]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b0000000011111111;
    wire [3:0] lut_436_select = {
                             in_data[158],
                             in_data[436],
                             in_data[751],
                             in_data[587]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b0001000100000001;
    wire [3:0] lut_437_select = {
                             in_data[200],
                             in_data[756],
                             in_data[690],
                             in_data[104]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b1110111011101110;
    wire [3:0] lut_438_select = {
                             in_data[728],
                             in_data[493],
                             in_data[543],
                             in_data[770]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b1110111111101111;
    wire [3:0] lut_439_select = {
                             in_data[763],
                             in_data[456],
                             in_data[772],
                             in_data[337]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b0001000000010000;
    wire [3:0] lut_440_select = {
                             in_data[281],
                             in_data[210],
                             in_data[740],
                             in_data[483]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b0010000000110000;
    wire [3:0] lut_441_select = {
                             in_data[534],
                             in_data[513],
                             in_data[693],
                             in_data[246]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b0011001100110011;
    wire [3:0] lut_442_select = {
                             in_data[725],
                             in_data[379],
                             in_data[631],
                             in_data[672]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1110111011111111;
    wire [3:0] lut_443_select = {
                             in_data[466],
                             in_data[783],
                             in_data[300],
                             in_data[105]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b1111000011110000;
    wire [3:0] lut_444_select = {
                             in_data[91],
                             in_data[329],
                             in_data[616],
                             in_data[716]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b1100111100001111;
    wire [3:0] lut_445_select = {
                             in_data[130],
                             in_data[544],
                             in_data[401],
                             in_data[57]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b0000010001010101;
    wire [3:0] lut_446_select = {
                             in_data[634],
                             in_data[776],
                             in_data[426],
                             in_data[637]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b1100110011101110;
    wire [3:0] lut_447_select = {
                             in_data[221],
                             in_data[319],
                             in_data[358],
                             in_data[489]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b0011001100110011;
    wire [3:0] lut_448_select = {
                             in_data[41],
                             in_data[602],
                             in_data[371],
                             in_data[564]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b0000111111001100;
    wire [3:0] lut_449_select = {
                             in_data[174],
                             in_data[169],
                             in_data[327],
                             in_data[700]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b1110111011101110;
    wire [3:0] lut_450_select = {
                             in_data[732],
                             in_data[639],
                             in_data[314],
                             in_data[579]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b0010001000110011;
    wire [3:0] lut_451_select = {
                             in_data[129],
                             in_data[87],
                             in_data[248],
                             in_data[367]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b0101000001010101;
    wire [3:0] lut_452_select = {
                             in_data[255],
                             in_data[667],
                             in_data[663],
                             in_data[175]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b0010101100000011;
    wire [3:0] lut_453_select = {
                             in_data[363],
                             in_data[469],
                             in_data[423],
                             in_data[254]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0000000000000011;
    wire [3:0] lut_454_select = {
                             in_data[435],
                             in_data[75],
                             in_data[65],
                             in_data[680]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b0000000011011101;
    wire [3:0] lut_455_select = {
                             in_data[274],
                             in_data[107],
                             in_data[650],
                             in_data[598]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b1111111111101110;
    wire [3:0] lut_456_select = {
                             in_data[465],
                             in_data[702],
                             in_data[712],
                             in_data[717]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b1111101011111010;
    wire [3:0] lut_457_select = {
                             in_data[590],
                             in_data[385],
                             in_data[173],
                             in_data[492]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b0101000011110000;
    wire [3:0] lut_458_select = {
                             in_data[256],
                             in_data[245],
                             in_data[141],
                             in_data[318]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b1111111100001100;
    wire [3:0] lut_459_select = {
                             in_data[275],
                             in_data[530],
                             in_data[233],
                             in_data[134]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b1011101010111010;
    wire [3:0] lut_460_select = {
                             in_data[699],
                             in_data[207],
                             in_data[143],
                             in_data[339]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b0100010001000100;
    wire [3:0] lut_461_select = {
                             in_data[168],
                             in_data[196],
                             in_data[409],
                             in_data[647]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b1111000011110011;
    wire [3:0] lut_462_select = {
                             in_data[38],
                             in_data[450],
                             in_data[538],
                             in_data[30]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b0000010101000111;
    wire [3:0] lut_463_select = {
                             in_data[360],
                             in_data[263],
                             in_data[425],
                             in_data[443]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b1100111111001111;
    wire [3:0] lut_464_select = {
                             in_data[671],
                             in_data[655],
                             in_data[80],
                             in_data[197]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b0100010100000000;
    wire [3:0] lut_465_select = {
                             in_data[292],
                             in_data[414],
                             in_data[595],
                             in_data[122]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b0000010011001100;
    wire [3:0] lut_466_select = {
                             in_data[573],
                             in_data[50],
                             in_data[262],
                             in_data[282]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1110110010101010;
    wire [3:0] lut_467_select = {
                             in_data[148],
                             in_data[726],
                             in_data[286],
                             in_data[345]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b0000001100000011;
    wire [3:0] lut_468_select = {
                             in_data[342],
                             in_data[623],
                             in_data[160],
                             in_data[63]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b1100111100000000;
    wire [3:0] lut_469_select = {
                             in_data[572],
                             in_data[390],
                             in_data[575],
                             in_data[109]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b0011000100110011;
    wire [3:0] lut_470_select = {
                             in_data[488],
                             in_data[480],
                             in_data[408],
                             in_data[696]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b1111111100110011;
    wire [3:0] lut_471_select = {
                             in_data[157],
                             in_data[28],
                             in_data[236],
                             in_data[420]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b0000110011001110;
    wire [3:0] lut_472_select = {
                             in_data[706],
                             in_data[668],
                             in_data[537],
                             in_data[540]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b0000000000000001;
    wire [3:0] lut_473_select = {
                             in_data[3],
                             in_data[536],
                             in_data[777],
                             in_data[172]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b0010000011110001;
    wire [3:0] lut_474_select = {
                             in_data[298],
                             in_data[288],
                             in_data[550],
                             in_data[524]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b1111111111101110;
    wire [3:0] lut_475_select = {
                             in_data[764],
                             in_data[120],
                             in_data[447],
                             in_data[266]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b0000000000000001;
    wire [3:0] lut_476_select = {
                             in_data[1],
                             in_data[82],
                             in_data[692],
                             in_data[424]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b1010101010101010;
    wire [3:0] lut_477_select = {
                             in_data[758],
                             in_data[39],
                             in_data[45],
                             in_data[624]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b0000000000000011;
    wire [3:0] lut_478_select = {
                             in_data[97],
                             in_data[392],
                             in_data[167],
                             in_data[4]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b1111101111111011;
    wire [3:0] lut_479_select = {
                             in_data[588],
                             in_data[226],
                             in_data[434],
                             in_data[558]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b1110101011101110;
    wire [3:0] lut_480_select = {
                             in_data[116],
                             in_data[496],
                             in_data[156],
                             in_data[215]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b0000111100001111;
    wire [3:0] lut_481_select = {
                             in_data[467],
                             in_data[268],
                             in_data[694],
                             in_data[60]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b1100110011001100;
    wire [3:0] lut_482_select = {
                             in_data[265],
                             in_data[526],
                             in_data[271],
                             in_data[346]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b0101010101010101;
    wire [3:0] lut_483_select = {
                             in_data[653],
                             in_data[611],
                             in_data[449],
                             in_data[713]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b0101010101010000;
    wire [3:0] lut_484_select = {
                             in_data[201],
                             in_data[159],
                             in_data[279],
                             in_data[151]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b0000000000000101;
    wire [3:0] lut_485_select = {
                             in_data[126],
                             in_data[439],
                             in_data[642],
                             in_data[94]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b0000111111000000;
    wire [3:0] lut_486_select = {
                             in_data[209],
                             in_data[330],
                             in_data[591],
                             in_data[51]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b1111110011111100;
    wire [3:0] lut_487_select = {
                             in_data[780],
                             in_data[528],
                             in_data[762],
                             in_data[56]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1010111110101010;
    wire [3:0] lut_488_select = {
                             in_data[70],
                             in_data[472],
                             in_data[646],
                             in_data[552]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b1100110011001101;
    wire [3:0] lut_489_select = {
                             in_data[22],
                             in_data[23],
                             in_data[675],
                             in_data[560]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b0000000000110010;
    wire [3:0] lut_490_select = {
                             in_data[164],
                             in_data[619],
                             in_data[208],
                             in_data[213]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b1111111100100010;
    wire [3:0] lut_491_select = {
                             in_data[242],
                             in_data[90],
                             in_data[546],
                             in_data[739]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b0000000000110011;
    wire [3:0] lut_492_select = {
                             in_data[412],
                             in_data[55],
                             in_data[441],
                             in_data[729]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b1111110111111101;
    wire [3:0] lut_493_select = {
                             in_data[62],
                             in_data[278],
                             in_data[387],
                             in_data[297]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b0010101001000101;
    wire [3:0] lut_494_select = {
                             in_data[267],
                             in_data[361],
                             in_data[497],
                             in_data[216]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b0000000001000100;
    wire [3:0] lut_495_select = {
                             in_data[498],
                             in_data[731],
                             in_data[461],
                             in_data[691]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b1111010111110101;
    wire [3:0] lut_496_select = {
                             in_data[505],
                             in_data[13],
                             in_data[24],
                             in_data[351]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b1111111110001001;
    wire [3:0] lut_497_select = {
                             in_data[135],
                             in_data[188],
                             in_data[484],
                             in_data[452]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b1111111111111100;
    wire [3:0] lut_498_select = {
                             in_data[306],
                             in_data[612],
                             in_data[253],
                             in_data[760]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b1111111111110000;
    wire [3:0] lut_499_select = {
                             in_data[499],
                             in_data[161],
                             in_data[648],
                             in_data[6]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b1010101010101011;
    wire [3:0] lut_500_select = {
                             in_data[451],
                             in_data[545],
                             in_data[198],
                             in_data[596]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b1110111110101110;
    wire [3:0] lut_501_select = {
                             in_data[765],
                             in_data[607],
                             in_data[437],
                             in_data[736]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b0101000000000010;
    wire [3:0] lut_502_select = {
                             in_data[608],
                             in_data[147],
                             in_data[260],
                             in_data[322]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b1111111110100000;
    wire [3:0] lut_503_select = {
                             in_data[659],
                             in_data[459],
                             in_data[117],
                             in_data[185]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b1011111110001010;
    wire [3:0] lut_504_select = {
                             in_data[603],
                             in_data[613],
                             in_data[471],
                             in_data[576]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b1111111111101110;
    wire [3:0] lut_505_select = {
                             in_data[626],
                             in_data[697],
                             in_data[710],
                             in_data[163]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b0011000100010001;
    wire [3:0] lut_506_select = {
                             in_data[133],
                             in_data[184],
                             in_data[368],
                             in_data[269]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b0000000000000001;
    wire [3:0] lut_507_select = {
                             in_data[140],
                             in_data[284],
                             in_data[741],
                             in_data[139]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b0000000000000001;
    wire [3:0] lut_508_select = {
                             in_data[309],
                             in_data[386],
                             in_data[714],
                             in_data[289]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b0001011101010000;
    wire [3:0] lut_509_select = {
                             in_data[688],
                             in_data[686],
                             in_data[584],
                             in_data[153]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b0000000000000001;
    wire [3:0] lut_510_select = {
                             in_data[81],
                             in_data[495],
                             in_data[78],
                             in_data[554]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0000000100000001;
    wire [3:0] lut_511_select = {
                             in_data[617],
                             in_data[604],
                             in_data[606],
                             in_data[333]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [15:0] lut_512_table = 16'b1101010111011100;
    wire [3:0] lut_512_select = {
                             in_data[561],
                             in_data[677],
                             in_data[556],
                             in_data[225]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [15:0] lut_513_table = 16'b1010111110101111;
    wire [3:0] lut_513_select = {
                             in_data[585],
                             in_data[464],
                             in_data[343],
                             in_data[750]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [15:0] lut_514_table = 16'b1110111111101111;
    wire [3:0] lut_514_select = {
                             in_data[76],
                             in_data[211],
                             in_data[400],
                             in_data[553]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [15:0] lut_515_table = 16'b1110101011101010;
    wire [3:0] lut_515_select = {
                             in_data[54],
                             in_data[67],
                             in_data[340],
                             in_data[239]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [15:0] lut_516_table = 16'b0000001100000000;
    wire [3:0] lut_516_select = {
                             in_data[516],
                             in_data[398],
                             in_data[506],
                             in_data[7]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [15:0] lut_517_table = 16'b1111110011111100;
    wire [3:0] lut_517_select = {
                             in_data[34],
                             in_data[721],
                             in_data[187],
                             in_data[391]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [15:0] lut_518_table = 16'b1111110011111100;
    wire [3:0] lut_518_select = {
                             in_data[673],
                             in_data[574],
                             in_data[231],
                             in_data[280]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [15:0] lut_519_table = 16'b0000001111110000;
    wire [3:0] lut_519_select = {
                             in_data[259],
                             in_data[214],
                             in_data[599],
                             in_data[406]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [15:0] lut_520_table = 16'b1010101110101010;
    wire [3:0] lut_520_select = {
                             in_data[517],
                             in_data[19],
                             in_data[562],
                             in_data[103]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [15:0] lut_521_table = 16'b1111111100000011;
    wire [3:0] lut_521_select = {
                             in_data[382],
                             in_data[630],
                             in_data[411],
                             in_data[338]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [15:0] lut_522_table = 16'b1111001111110011;
    wire [3:0] lut_522_select = {
                             in_data[224],
                             in_data[567],
                             in_data[237],
                             in_data[21]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [15:0] lut_523_table = 16'b0000000011111111;
    wire [3:0] lut_523_select = {
                             in_data[244],
                             in_data[479],
                             in_data[194],
                             in_data[113]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [15:0] lut_524_table = 16'b0000000100000001;
    wire [3:0] lut_524_select = {
                             in_data[85],
                             in_data[15],
                             in_data[635],
                             in_data[114]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [15:0] lut_525_table = 16'b1000010110100101;
    wire [3:0] lut_525_select = {
                             in_data[36],
                             in_data[186],
                             in_data[405],
                             in_data[628]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [15:0] lut_526_table = 16'b0100000101000011;
    wire [3:0] lut_526_select = {
                             in_data[42],
                             in_data[326],
                             in_data[388],
                             in_data[369]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [15:0] lut_527_table = 16'b0001000100000000;
    wire [3:0] lut_527_select = {
                             in_data[404],
                             in_data[335],
                             in_data[74],
                             in_data[622]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [15:0] lut_528_table = 16'b0010111100100010;
    wire [3:0] lut_528_select = {
                             in_data[518],
                             in_data[121],
                             in_data[600],
                             in_data[227]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [15:0] lut_529_table = 16'b0000111100001111;
    wire [3:0] lut_529_select = {
                             in_data[308],
                             in_data[597],
                             in_data[191],
                             in_data[615]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [15:0] lut_530_table = 16'b1111000011110001;
    wire [3:0] lut_530_select = {
                             in_data[132],
                             in_data[359],
                             in_data[504],
                             in_data[416]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [15:0] lut_531_table = 16'b0000111100001111;
    wire [3:0] lut_531_select = {
                             in_data[199],
                             in_data[548],
                             in_data[722],
                             in_data[136]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [15:0] lut_532_table = 16'b1110111111001100;
    wire [3:0] lut_532_select = {
                             in_data[601],
                             in_data[718],
                             in_data[101],
                             in_data[440]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [15:0] lut_533_table = 16'b1111111111110011;
    wire [3:0] lut_533_select = {
                             in_data[35],
                             in_data[641],
                             in_data[559],
                             in_data[53]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [15:0] lut_534_table = 16'b1110100011111110;
    wire [3:0] lut_534_select = {
                             in_data[312],
                             in_data[670],
                             in_data[73],
                             in_data[44]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [15:0] lut_535_table = 16'b1111010001111110;
    wire [3:0] lut_535_select = {
                             in_data[234],
                             in_data[182],
                             in_data[93],
                             in_data[240]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [15:0] lut_536_table = 16'b0000011100001111;
    wire [3:0] lut_536_select = {
                             in_data[238],
                             in_data[377],
                             in_data[511],
                             in_data[145]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [15:0] lut_537_table = 16'b0000000011111100;
    wire [3:0] lut_537_select = {
                             in_data[470],
                             in_data[321],
                             in_data[715],
                             in_data[487]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [15:0] lut_538_table = 16'b1100000011110011;
    wire [3:0] lut_538_select = {
                             in_data[313],
                             in_data[719],
                             in_data[232],
                             in_data[27]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [15:0] lut_539_table = 16'b0000110000001111;
    wire [3:0] lut_539_select = {
                             in_data[551],
                             in_data[108],
                             in_data[689],
                             in_data[52]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [15:0] lut_540_table = 16'b1111000011110000;
    wire [3:0] lut_540_select = {
                             in_data[395],
                             in_data[311],
                             in_data[759],
                             in_data[421]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [15:0] lut_541_table = 16'b1100110011101110;
    wire [3:0] lut_541_select = {
                             in_data[746],
                             in_data[365],
                             in_data[743],
                             in_data[491]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [15:0] lut_542_table = 16'b1111111111110101;
    wire [3:0] lut_542_select = {
                             in_data[79],
                             in_data[247],
                             in_data[110],
                             in_data[241]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [15:0] lut_543_table = 16'b0100010001010101;
    wire [3:0] lut_543_select = {
                             in_data[328],
                             in_data[12],
                             in_data[389],
                             in_data[190]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [15:0] lut_544_table = 16'b1111111111111100;
    wire [3:0] lut_544_select = {
                             in_data[705],
                             in_data[769],
                             in_data[294],
                             in_data[482]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [15:0] lut_545_table = 16'b1111111111111000;
    wire [3:0] lut_545_select = {
                             in_data[296],
                             in_data[98],
                             in_data[325],
                             in_data[651]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [15:0] lut_546_table = 16'b0011111111110000;
    wire [3:0] lut_546_select = {
                             in_data[625],
                             in_data[656],
                             in_data[258],
                             in_data[222]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [15:0] lut_547_table = 16'b0000010100000001;
    wire [3:0] lut_547_select = {
                             in_data[766],
                             in_data[102],
                             in_data[781],
                             in_data[666]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [15:0] lut_548_table = 16'b0100010100000101;
    wire [3:0] lut_548_select = {
                             in_data[307],
                             in_data[431],
                             in_data[177],
                             in_data[514]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [15:0] lut_549_table = 16'b1111111111110000;
    wire [3:0] lut_549_select = {
                             in_data[563],
                             in_data[711],
                             in_data[112],
                             in_data[166]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [15:0] lut_550_table = 16'b0000000100000001;
    wire [3:0] lut_550_select = {
                             in_data[753],
                             in_data[761],
                             in_data[202],
                             in_data[228]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [15:0] lut_551_table = 16'b0000111100001111;
    wire [3:0] lut_551_select = {
                             in_data[709],
                             in_data[181],
                             in_data[86],
                             in_data[727]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [15:0] lut_552_table = 16'b1101110101000101;
    wire [3:0] lut_552_select = {
                             in_data[748],
                             in_data[204],
                             in_data[723],
                             in_data[118]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [15:0] lut_553_table = 16'b1111110000001100;
    wire [3:0] lut_553_select = {
                             in_data[127],
                             in_data[95],
                             in_data[295],
                             in_data[384]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [15:0] lut_554_table = 16'b1111111111001111;
    wire [3:0] lut_554_select = {
                             in_data[557],
                             in_data[374],
                             in_data[582],
                             in_data[20]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [15:0] lut_555_table = 16'b1111000011111111;
    wire [3:0] lut_555_select = {
                             in_data[533],
                             in_data[720],
                             in_data[643],
                             in_data[49]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [15:0] lut_556_table = 16'b1111111111101110;
    wire [3:0] lut_556_select = {
                             in_data[678],
                             in_data[170],
                             in_data[468],
                             in_data[509]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [15:0] lut_557_table = 16'b0111001101110011;
    wire [3:0] lut_557_select = {
                             in_data[46],
                             in_data[654],
                             in_data[235],
                             in_data[383]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [15:0] lut_558_table = 16'b0000000010101010;
    wire [3:0] lut_558_select = {
                             in_data[512],
                             in_data[84],
                             in_data[448],
                             in_data[264]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [15:0] lut_559_table = 16'b0000000000000001;
    wire [3:0] lut_559_select = {
                             in_data[138],
                             in_data[33],
                             in_data[303],
                             in_data[738]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [15:0] lut_560_table = 16'b1111111110101010;
    wire [3:0] lut_560_select = {
                             in_data[331],
                             in_data[757],
                             in_data[679],
                             in_data[273]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [15:0] lut_561_table = 16'b0001000100010001;
    wire [3:0] lut_561_select = {
                             in_data[394],
                             in_data[315],
                             in_data[96],
                             in_data[149]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [15:0] lut_562_table = 16'b1111111111111110;
    wire [3:0] lut_562_select = {
                             in_data[37],
                             in_data[100],
                             in_data[737],
                             in_data[61]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [15:0] lut_563_table = 16'b1101110011011100;
    wire [3:0] lut_563_select = {
                             in_data[58],
                             in_data[586],
                             in_data[541],
                             in_data[287]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [15:0] lut_564_table = 16'b0101000011110101;
    wire [3:0] lut_564_select = {
                             in_data[707],
                             in_data[510],
                             in_data[83],
                             in_data[380]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [15:0] lut_565_table = 16'b0010111110101111;
    wire [3:0] lut_565_select = {
                             in_data[477],
                             in_data[270],
                             in_data[355],
                             in_data[376]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [15:0] lut_566_table = 16'b1111111111001100;
    wire [3:0] lut_566_select = {
                             in_data[399],
                             in_data[645],
                             in_data[347],
                             in_data[486]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [15:0] lut_567_table = 16'b0000000000000011;
    wire [3:0] lut_567_select = {
                             in_data[131],
                             in_data[539],
                             in_data[119],
                             in_data[520]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [15:0] lut_568_table = 16'b0000000000110011;
    wire [3:0] lut_568_select = {
                             in_data[128],
                             in_data[755],
                             in_data[633],
                             in_data[88]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [15:0] lut_569_table = 16'b1110110011111110;
    wire [3:0] lut_569_select = {
                             in_data[301],
                             in_data[669],
                             in_data[155],
                             in_data[500]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [15:0] lut_570_table = 16'b0000000000010001;
    wire [3:0] lut_570_select = {
                             in_data[125],
                             in_data[703],
                             in_data[583],
                             in_data[507]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [15:0] lut_571_table = 16'b1010101010100010;
    wire [3:0] lut_571_select = {
                             in_data[261],
                             in_data[660],
                             in_data[508],
                             in_data[373]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [15:0] lut_572_table = 16'b1111111101010101;
    wire [3:0] lut_572_select = {
                             in_data[593],
                             in_data[614],
                             in_data[531],
                             in_data[344]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [15:0] lut_573_table = 16'b1111111100000100;
    wire [3:0] lut_573_select = {
                             in_data[357],
                             in_data[162],
                             in_data[519],
                             in_data[48]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [15:0] lut_574_table = 16'b1010000011111010;
    wire [3:0] lut_574_select = {
                             in_data[733],
                             in_data[40],
                             in_data[754],
                             in_data[768]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [15:0] lut_575_table = 16'b1111000111110001;
    wire [3:0] lut_575_select = {
                             in_data[336],
                             in_data[66],
                             in_data[299],
                             in_data[775]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [15:0] lut_576_table = 16'b0011001000110011;
    wire [3:0] lut_576_select = {
                             in_data[77],
                             in_data[620],
                             in_data[485],
                             in_data[724]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [15:0] lut_577_table = 16'b0101000001010000;
    wire [3:0] lut_577_select = {
                             in_data[144],
                             in_data[350],
                             in_data[503],
                             in_data[501]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [15:0] lut_578_table = 16'b1110111011101110;
    wire [3:0] lut_578_select = {
                             in_data[419],
                             in_data[16],
                             in_data[636],
                             in_data[410]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [15:0] lut_579_table = 16'b1111111101010101;
    wire [3:0] lut_579_select = {
                             in_data[577],
                             in_data[478],
                             in_data[393],
                             in_data[460]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [15:0] lut_580_table = 16'b1111111011110101;
    wire [3:0] lut_580_select = {
                             in_data[353],
                             in_data[522],
                             in_data[68],
                             in_data[462]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [15:0] lut_581_table = 16'b0000000000000001;
    wire [3:0] lut_581_select = {
                             in_data[446],
                             in_data[277],
                             in_data[43],
                             in_data[29]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [15:0] lut_582_table = 16'b1111000111110011;
    wire [3:0] lut_582_select = {
                             in_data[217],
                             in_data[415],
                             in_data[378],
                             in_data[150]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [15:0] lut_583_table = 16'b0000111100001100;
    wire [3:0] lut_583_select = {
                             in_data[767],
                             in_data[332],
                             in_data[205],
                             in_data[2]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [15:0] lut_584_table = 16'b0000111101001111;
    wire [3:0] lut_584_select = {
                             in_data[683],
                             in_data[515],
                             in_data[749],
                             in_data[527]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [15:0] lut_585_table = 16'b0100010001001100;
    wire [3:0] lut_585_select = {
                             in_data[251],
                             in_data[589],
                             in_data[565],
                             in_data[89]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [15:0] lut_586_table = 16'b1111111101001100;
    wire [3:0] lut_586_select = {
                             in_data[581],
                             in_data[5],
                             in_data[0],
                             in_data[111]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [15:0] lut_587_table = 16'b1111011101110000;
    wire [3:0] lut_587_select = {
                             in_data[366],
                             in_data[555],
                             in_data[674],
                             in_data[532]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [15:0] lut_588_table = 16'b1010010000000101;
    wire [3:0] lut_588_select = {
                             in_data[179],
                             in_data[150],
                             in_data[562],
                             in_data[372]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [15:0] lut_589_table = 16'b0000001100000011;
    wire [3:0] lut_589_select = {
                             in_data[55],
                             in_data[247],
                             in_data[358],
                             in_data[3]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [15:0] lut_590_table = 16'b0000000000001010;
    wire [3:0] lut_590_select = {
                             in_data[430],
                             in_data[455],
                             in_data[13],
                             in_data[407]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [15:0] lut_591_table = 16'b1111111111110010;
    wire [3:0] lut_591_select = {
                             in_data[92],
                             in_data[460],
                             in_data[627],
                             in_data[104]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [15:0] lut_592_table = 16'b1110110011111000;
    wire [3:0] lut_592_select = {
                             in_data[345],
                             in_data[690],
                             in_data[491],
                             in_data[327]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [15:0] lut_593_table = 16'b1100000011111100;
    wire [3:0] lut_593_select = {
                             in_data[251],
                             in_data[602],
                             in_data[474],
                             in_data[589]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [15:0] lut_594_table = 16'b0010101010101011;
    wire [3:0] lut_594_select = {
                             in_data[531],
                             in_data[635],
                             in_data[419],
                             in_data[739]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [15:0] lut_595_table = 16'b0001000000010000;
    wire [3:0] lut_595_select = {
                             in_data[84],
                             in_data[27],
                             in_data[48],
                             in_data[166]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [15:0] lut_596_table = 16'b0000000100000001;
    wire [3:0] lut_596_select = {
                             in_data[146],
                             in_data[383],
                             in_data[457],
                             in_data[96]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [15:0] lut_597_table = 16'b0000111100101010;
    wire [3:0] lut_597_select = {
                             in_data[303],
                             in_data[444],
                             in_data[62],
                             in_data[367]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [15:0] lut_598_table = 16'b0000000000010101;
    wire [3:0] lut_598_select = {
                             in_data[441],
                             in_data[773],
                             in_data[713],
                             in_data[735]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [15:0] lut_599_table = 16'b0100110011001100;
    wire [3:0] lut_599_select = {
                             in_data[40],
                             in_data[400],
                             in_data[624],
                             in_data[102]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [15:0] lut_600_table = 16'b1111101111111011;
    wire [3:0] lut_600_select = {
                             in_data[716],
                             in_data[98],
                             in_data[287],
                             in_data[745]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [15:0] lut_601_table = 16'b1111111111110000;
    wire [3:0] lut_601_select = {
                             in_data[640],
                             in_data[245],
                             in_data[705],
                             in_data[533]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [15:0] lut_602_table = 16'b1111111111111100;
    wire [3:0] lut_602_select = {
                             in_data[329],
                             in_data[743],
                             in_data[357],
                             in_data[698]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [15:0] lut_603_table = 16'b0000011100000001;
    wire [3:0] lut_603_select = {
                             in_data[119],
                             in_data[191],
                             in_data[223],
                             in_data[132]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [15:0] lut_604_table = 16'b0000000100000011;
    wire [3:0] lut_604_select = {
                             in_data[23],
                             in_data[579],
                             in_data[494],
                             in_data[769]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [15:0] lut_605_table = 16'b0000110011001110;
    wire [3:0] lut_605_select = {
                             in_data[408],
                             in_data[74],
                             in_data[355],
                             in_data[285]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [15:0] lut_606_table = 16'b1111111100001101;
    wire [3:0] lut_606_select = {
                             in_data[272],
                             in_data[451],
                             in_data[228],
                             in_data[325]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [15:0] lut_607_table = 16'b1111111111101111;
    wire [3:0] lut_607_select = {
                             in_data[222],
                             in_data[435],
                             in_data[44],
                             in_data[535]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [15:0] lut_608_table = 16'b0000000010101011;
    wire [3:0] lut_608_select = {
                             in_data[260],
                             in_data[61],
                             in_data[761],
                             in_data[254]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [15:0] lut_609_table = 16'b0000000000110011;
    wire [3:0] lut_609_select = {
                             in_data[155],
                             in_data[449],
                             in_data[344],
                             in_data[561]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [15:0] lut_610_table = 16'b0000101000001010;
    wire [3:0] lut_610_select = {
                             in_data[35],
                             in_data[507],
                             in_data[11],
                             in_data[543]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [15:0] lut_611_table = 16'b0000010000000101;
    wire [3:0] lut_611_select = {
                             in_data[316],
                             in_data[481],
                             in_data[168],
                             in_data[232]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [15:0] lut_612_table = 16'b0000010001000101;
    wire [3:0] lut_612_select = {
                             in_data[115],
                             in_data[42],
                             in_data[334],
                             in_data[704]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [15:0] lut_613_table = 16'b1111111110101010;
    wire [3:0] lut_613_select = {
                             in_data[508],
                             in_data[614],
                             in_data[43],
                             in_data[497]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [15:0] lut_614_table = 16'b1011001111110011;
    wire [3:0] lut_614_select = {
                             in_data[674],
                             in_data[127],
                             in_data[404],
                             in_data[53]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [15:0] lut_615_table = 16'b0000111100001111;
    wire [3:0] lut_615_select = {
                             in_data[346],
                             in_data[515],
                             in_data[10],
                             in_data[341]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [15:0] lut_616_table = 16'b1111111101010101;
    wire [3:0] lut_616_select = {
                             in_data[485],
                             in_data[439],
                             in_data[418],
                             in_data[207]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [15:0] lut_617_table = 16'b1111010111110000;
    wire [3:0] lut_617_select = {
                             in_data[566],
                             in_data[378],
                             in_data[724],
                             in_data[261]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [15:0] lut_618_table = 16'b1010101110101010;
    wire [3:0] lut_618_select = {
                             in_data[524],
                             in_data[767],
                             in_data[388],
                             in_data[186]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [15:0] lut_619_table = 16'b1011101010101010;
    wire [3:0] lut_619_select = {
                             in_data[764],
                             in_data[634],
                             in_data[527],
                             in_data[213]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [15:0] lut_620_table = 16'b1010000011110000;
    wire [3:0] lut_620_select = {
                             in_data[734],
                             in_data[348],
                             in_data[783],
                             in_data[663]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [15:0] lut_621_table = 16'b1111000011111111;
    wire [3:0] lut_621_select = {
                             in_data[630],
                             in_data[513],
                             in_data[392],
                             in_data[90]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [15:0] lut_622_table = 16'b0000111100000011;
    wire [3:0] lut_622_select = {
                             in_data[205],
                             in_data[453],
                             in_data[187],
                             in_data[22]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [15:0] lut_623_table = 16'b1111001111111011;
    wire [3:0] lut_623_select = {
                             in_data[462],
                             in_data[152],
                             in_data[296],
                             in_data[163]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [15:0] lut_624_table = 16'b1010101110101011;
    wire [3:0] lut_624_select = {
                             in_data[417],
                             in_data[249],
                             in_data[521],
                             in_data[414]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [15:0] lut_625_table = 16'b1111111111110000;
    wire [3:0] lut_625_select = {
                             in_data[737],
                             in_data[204],
                             in_data[148],
                             in_data[25]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [15:0] lut_626_table = 16'b0011001100110011;
    wire [3:0] lut_626_select = {
                             in_data[520],
                             in_data[505],
                             in_data[184],
                             in_data[756]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [15:0] lut_627_table = 16'b0111011100010001;
    wire [3:0] lut_627_select = {
                             in_data[71],
                             in_data[749],
                             in_data[190],
                             in_data[248]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [15:0] lut_628_table = 16'b1111011101000000;
    wire [3:0] lut_628_select = {
                             in_data[219],
                             in_data[525],
                             in_data[607],
                             in_data[512]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [15:0] lut_629_table = 16'b0011001100000000;
    wire [3:0] lut_629_select = {
                             in_data[265],
                             in_data[24],
                             in_data[151],
                             in_data[565]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [15:0] lut_630_table = 16'b0000000011001100;
    wire [3:0] lut_630_select = {
                             in_data[661],
                             in_data[598],
                             in_data[459],
                             in_data[727]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [15:0] lut_631_table = 16'b1011101010110000;
    wire [3:0] lut_631_select = {
                             in_data[465],
                             in_data[244],
                             in_data[109],
                             in_data[658]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [15:0] lut_632_table = 16'b0101111100001111;
    wire [3:0] lut_632_select = {
                             in_data[311],
                             in_data[351],
                             in_data[385],
                             in_data[125]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [15:0] lut_633_table = 16'b1111111011111010;
    wire [3:0] lut_633_select = {
                             in_data[567],
                             in_data[188],
                             in_data[645],
                             in_data[662]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [15:0] lut_634_table = 16'b0000000000100010;
    wire [3:0] lut_634_select = {
                             in_data[592],
                             in_data[169],
                             in_data[94],
                             in_data[270]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [15:0] lut_635_table = 16'b0101000101010101;
    wire [3:0] lut_635_select = {
                             in_data[708],
                             in_data[519],
                             in_data[568],
                             in_data[654]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [15:0] lut_636_table = 16'b0011000100010000;
    wire [3:0] lut_636_select = {
                             in_data[778],
                             in_data[320],
                             in_data[618],
                             in_data[726]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [15:0] lut_637_table = 16'b1110111011111111;
    wire [3:0] lut_637_select = {
                             in_data[603],
                             in_data[768],
                             in_data[637],
                             in_data[709]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [15:0] lut_638_table = 16'b0000111100001111;
    wire [3:0] lut_638_select = {
                             in_data[755],
                             in_data[381],
                             in_data[680],
                             in_data[777]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [15:0] lut_639_table = 16'b1100110011001111;
    wire [3:0] lut_639_select = {
                             in_data[625],
                             in_data[539],
                             in_data[176],
                             in_data[558]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
    
    // LUT : 640
    wire [15:0] lut_640_table = 16'b1111111110101010;
    wire [3:0] lut_640_select = {
                             in_data[511],
                             in_data[782],
                             in_data[677],
                             in_data[669]};
    
    wire lut_640_out = lut_640_table[lut_640_select];
    
    generate
    if ( USE_REG ) begin : ff_640
        reg   lut_640_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_640_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_640_ff <= lut_640_out;
            end
        end
        
        assign out_data[640] = lut_640_ff;
    end
    else begin : no_ff_640
        assign out_data[640] = lut_640_out;
    end
    endgenerate
    
    
    
    // LUT : 641
    wire [15:0] lut_641_table = 16'b1111111111110000;
    wire [3:0] lut_641_select = {
                             in_data[717],
                             in_data[409],
                             in_data[393],
                             in_data[17]};
    
    wire lut_641_out = lut_641_table[lut_641_select];
    
    generate
    if ( USE_REG ) begin : ff_641
        reg   lut_641_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_641_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_641_ff <= lut_641_out;
            end
        end
        
        assign out_data[641] = lut_641_ff;
    end
    else begin : no_ff_641
        assign out_data[641] = lut_641_out;
    end
    endgenerate
    
    
    
    // LUT : 642
    wire [15:0] lut_642_table = 16'b0011000000110011;
    wire [3:0] lut_642_select = {
                             in_data[319],
                             in_data[503],
                             in_data[38],
                             in_data[308]};
    
    wire lut_642_out = lut_642_table[lut_642_select];
    
    generate
    if ( USE_REG ) begin : ff_642
        reg   lut_642_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_642_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_642_ff <= lut_642_out;
            end
        end
        
        assign out_data[642] = lut_642_ff;
    end
    else begin : no_ff_642
        assign out_data[642] = lut_642_out;
    end
    endgenerate
    
    
    
    // LUT : 643
    wire [15:0] lut_643_table = 16'b0011001100110011;
    wire [3:0] lut_643_select = {
                             in_data[696],
                             in_data[751],
                             in_data[571],
                             in_data[534]};
    
    wire lut_643_out = lut_643_table[lut_643_select];
    
    generate
    if ( USE_REG ) begin : ff_643
        reg   lut_643_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_643_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_643_ff <= lut_643_out;
            end
        end
        
        assign out_data[643] = lut_643_ff;
    end
    else begin : no_ff_643
        assign out_data[643] = lut_643_out;
    end
    endgenerate
    
    
    
    // LUT : 644
    wire [15:0] lut_644_table = 16'b1011101010111010;
    wire [3:0] lut_644_select = {
                             in_data[39],
                             in_data[280],
                             in_data[468],
                             in_data[538]};
    
    wire lut_644_out = lut_644_table[lut_644_select];
    
    generate
    if ( USE_REG ) begin : ff_644
        reg   lut_644_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_644_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_644_ff <= lut_644_out;
            end
        end
        
        assign out_data[644] = lut_644_ff;
    end
    else begin : no_ff_644
        assign out_data[644] = lut_644_out;
    end
    endgenerate
    
    
    
    // LUT : 645
    wire [15:0] lut_645_table = 16'b0000000011001100;
    wire [3:0] lut_645_select = {
                             in_data[694],
                             in_data[229],
                             in_data[629],
                             in_data[328]};
    
    wire lut_645_out = lut_645_table[lut_645_select];
    
    generate
    if ( USE_REG ) begin : ff_645
        reg   lut_645_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_645_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_645_ff <= lut_645_out;
            end
        end
        
        assign out_data[645] = lut_645_ff;
    end
    else begin : no_ff_645
        assign out_data[645] = lut_645_out;
    end
    endgenerate
    
    
    
    // LUT : 646
    wire [15:0] lut_646_table = 16'b0011000000110011;
    wire [3:0] lut_646_select = {
                             in_data[284],
                             in_data[500],
                             in_data[714],
                             in_data[336]};
    
    wire lut_646_out = lut_646_table[lut_646_select];
    
    generate
    if ( USE_REG ) begin : ff_646
        reg   lut_646_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_646_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_646_ff <= lut_646_out;
            end
        end
        
        assign out_data[646] = lut_646_ff;
    end
    else begin : no_ff_646
        assign out_data[646] = lut_646_out;
    end
    endgenerate
    
    
    
    // LUT : 647
    wire [15:0] lut_647_table = 16'b1101111100010001;
    wire [3:0] lut_647_select = {
                             in_data[428],
                             in_data[12],
                             in_data[200],
                             in_data[597]};
    
    wire lut_647_out = lut_647_table[lut_647_select];
    
    generate
    if ( USE_REG ) begin : ff_647
        reg   lut_647_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_647_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_647_ff <= lut_647_out;
            end
        end
        
        assign out_data[647] = lut_647_ff;
    end
    else begin : no_ff_647
        assign out_data[647] = lut_647_out;
    end
    endgenerate
    
    
    
    // LUT : 648
    wire [15:0] lut_648_table = 16'b0100110011111110;
    wire [3:0] lut_648_select = {
                             in_data[161],
                             in_data[206],
                             in_data[128],
                             in_data[496]};
    
    wire lut_648_out = lut_648_table[lut_648_select];
    
    generate
    if ( USE_REG ) begin : ff_648
        reg   lut_648_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_648_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_648_ff <= lut_648_out;
            end
        end
        
        assign out_data[648] = lut_648_ff;
    end
    else begin : no_ff_648
        assign out_data[648] = lut_648_out;
    end
    endgenerate
    
    
    
    // LUT : 649
    wire [15:0] lut_649_table = 16'b1111111111111100;
    wire [3:0] lut_649_select = {
                             in_data[556],
                             in_data[154],
                             in_data[529],
                             in_data[208]};
    
    wire lut_649_out = lut_649_table[lut_649_select];
    
    generate
    if ( USE_REG ) begin : ff_649
        reg   lut_649_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_649_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_649_ff <= lut_649_out;
            end
        end
        
        assign out_data[649] = lut_649_ff;
    end
    else begin : no_ff_649
        assign out_data[649] = lut_649_out;
    end
    endgenerate
    
    
    
    // LUT : 650
    wire [15:0] lut_650_table = 16'b1111111110100010;
    wire [3:0] lut_650_select = {
                             in_data[670],
                             in_data[2],
                             in_data[617],
                             in_data[729]};
    
    wire lut_650_out = lut_650_table[lut_650_select];
    
    generate
    if ( USE_REG ) begin : ff_650
        reg   lut_650_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_650_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_650_ff <= lut_650_out;
            end
        end
        
        assign out_data[650] = lut_650_ff;
    end
    else begin : no_ff_650
        assign out_data[650] = lut_650_out;
    end
    endgenerate
    
    
    
    // LUT : 651
    wire [15:0] lut_651_table = 16'b0011001110110011;
    wire [3:0] lut_651_select = {
                             in_data[192],
                             in_data[332],
                             in_data[631],
                             in_data[81]};
    
    wire lut_651_out = lut_651_table[lut_651_select];
    
    generate
    if ( USE_REG ) begin : ff_651
        reg   lut_651_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_651_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_651_ff <= lut_651_out;
            end
        end
        
        assign out_data[651] = lut_651_ff;
    end
    else begin : no_ff_651
        assign out_data[651] = lut_651_out;
    end
    endgenerate
    
    
    
    // LUT : 652
    wire [15:0] lut_652_table = 16'b1111111111110000;
    wire [3:0] lut_652_select = {
                             in_data[246],
                             in_data[471],
                             in_data[195],
                             in_data[532]};
    
    wire lut_652_out = lut_652_table[lut_652_select];
    
    generate
    if ( USE_REG ) begin : ff_652
        reg   lut_652_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_652_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_652_ff <= lut_652_out;
            end
        end
        
        assign out_data[652] = lut_652_ff;
    end
    else begin : no_ff_652
        assign out_data[652] = lut_652_out;
    end
    endgenerate
    
    
    
    // LUT : 653
    wire [15:0] lut_653_table = 16'b1111111111001100;
    wire [3:0] lut_653_select = {
                             in_data[134],
                             in_data[215],
                             in_data[429],
                             in_data[7]};
    
    wire lut_653_out = lut_653_table[lut_653_select];
    
    generate
    if ( USE_REG ) begin : ff_653
        reg   lut_653_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_653_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_653_ff <= lut_653_out;
            end
        end
        
        assign out_data[653] = lut_653_ff;
    end
    else begin : no_ff_653
        assign out_data[653] = lut_653_out;
    end
    endgenerate
    
    
    
    // LUT : 654
    wire [15:0] lut_654_table = 16'b1111111110101011;
    wire [3:0] lut_654_select = {
                             in_data[374],
                             in_data[144],
                             in_data[211],
                             in_data[343]};
    
    wire lut_654_out = lut_654_table[lut_654_select];
    
    generate
    if ( USE_REG ) begin : ff_654
        reg   lut_654_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_654_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_654_ff <= lut_654_out;
            end
        end
        
        assign out_data[654] = lut_654_ff;
    end
    else begin : no_ff_654
        assign out_data[654] = lut_654_out;
    end
    endgenerate
    
    
    
    // LUT : 655
    wire [15:0] lut_655_table = 16'b0000000000100010;
    wire [3:0] lut_655_select = {
                             in_data[37],
                             in_data[29],
                             in_data[91],
                             in_data[557]};
    
    wire lut_655_out = lut_655_table[lut_655_select];
    
    generate
    if ( USE_REG ) begin : ff_655
        reg   lut_655_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_655_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_655_ff <= lut_655_out;
            end
        end
        
        assign out_data[655] = lut_655_ff;
    end
    else begin : no_ff_655
        assign out_data[655] = lut_655_out;
    end
    endgenerate
    
    
    
    // LUT : 656
    wire [15:0] lut_656_table = 16'b0101000101010001;
    wire [3:0] lut_656_select = {
                             in_data[421],
                             in_data[484],
                             in_data[445],
                             in_data[237]};
    
    wire lut_656_out = lut_656_table[lut_656_select];
    
    generate
    if ( USE_REG ) begin : ff_656
        reg   lut_656_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_656_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_656_ff <= lut_656_out;
            end
        end
        
        assign out_data[656] = lut_656_ff;
    end
    else begin : no_ff_656
        assign out_data[656] = lut_656_out;
    end
    endgenerate
    
    
    
    // LUT : 657
    wire [15:0] lut_657_table = 16'b0000001100000011;
    wire [3:0] lut_657_select = {
                             in_data[79],
                             in_data[578],
                             in_data[547],
                             in_data[49]};
    
    wire lut_657_out = lut_657_table[lut_657_select];
    
    generate
    if ( USE_REG ) begin : ff_657
        reg   lut_657_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_657_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_657_ff <= lut_657_out;
            end
        end
        
        assign out_data[657] = lut_657_ff;
    end
    else begin : no_ff_657
        assign out_data[657] = lut_657_out;
    end
    endgenerate
    
    
    
    // LUT : 658
    wire [15:0] lut_658_table = 16'b0001000001110101;
    wire [3:0] lut_658_select = {
                             in_data[549],
                             in_data[123],
                             in_data[456],
                             in_data[576]};
    
    wire lut_658_out = lut_658_table[lut_658_select];
    
    generate
    if ( USE_REG ) begin : ff_658
        reg   lut_658_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_658_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_658_ff <= lut_658_out;
            end
        end
        
        assign out_data[658] = lut_658_ff;
    end
    else begin : no_ff_658
        assign out_data[658] = lut_658_out;
    end
    endgenerate
    
    
    
    // LUT : 659
    wire [15:0] lut_659_table = 16'b1111111110111011;
    wire [3:0] lut_659_select = {
                             in_data[473],
                             in_data[28],
                             in_data[209],
                             in_data[638]};
    
    wire lut_659_out = lut_659_table[lut_659_select];
    
    generate
    if ( USE_REG ) begin : ff_659
        reg   lut_659_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_659_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_659_ff <= lut_659_out;
            end
        end
        
        assign out_data[659] = lut_659_ff;
    end
    else begin : no_ff_659
        assign out_data[659] = lut_659_out;
    end
    endgenerate
    
    
    
    // LUT : 660
    wire [15:0] lut_660_table = 16'b0011001100110011;
    wire [3:0] lut_660_select = {
                             in_data[315],
                             in_data[641],
                             in_data[509],
                             in_data[689]};
    
    wire lut_660_out = lut_660_table[lut_660_select];
    
    generate
    if ( USE_REG ) begin : ff_660
        reg   lut_660_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_660_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_660_ff <= lut_660_out;
            end
        end
        
        assign out_data[660] = lut_660_ff;
    end
    else begin : no_ff_660
        assign out_data[660] = lut_660_out;
    end
    endgenerate
    
    
    
    // LUT : 661
    wire [15:0] lut_661_table = 16'b1111000011111111;
    wire [3:0] lut_661_select = {
                             in_data[412],
                             in_data[707],
                             in_data[173],
                             in_data[781]};
    
    wire lut_661_out = lut_661_table[lut_661_select];
    
    generate
    if ( USE_REG ) begin : ff_661
        reg   lut_661_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_661_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_661_ff <= lut_661_out;
            end
        end
        
        assign out_data[661] = lut_661_ff;
    end
    else begin : no_ff_661
        assign out_data[661] = lut_661_out;
    end
    endgenerate
    
    
    
    // LUT : 662
    wire [15:0] lut_662_table = 16'b1111101011111010;
    wire [3:0] lut_662_select = {
                             in_data[85],
                             in_data[360],
                             in_data[8],
                             in_data[628]};
    
    wire lut_662_out = lut_662_table[lut_662_select];
    
    generate
    if ( USE_REG ) begin : ff_662
        reg   lut_662_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_662_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_662_ff <= lut_662_out;
            end
        end
        
        assign out_data[662] = lut_662_ff;
    end
    else begin : no_ff_662
        assign out_data[662] = lut_662_out;
    end
    endgenerate
    
    
    
    // LUT : 663
    wire [15:0] lut_663_table = 16'b0000101100001011;
    wire [3:0] lut_663_select = {
                             in_data[588],
                             in_data[427],
                             in_data[495],
                             in_data[770]};
    
    wire lut_663_out = lut_663_table[lut_663_select];
    
    generate
    if ( USE_REG ) begin : ff_663
        reg   lut_663_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_663_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_663_ff <= lut_663_out;
            end
        end
        
        assign out_data[663] = lut_663_ff;
    end
    else begin : no_ff_663
        assign out_data[663] = lut_663_out;
    end
    endgenerate
    
    
    
    // LUT : 664
    wire [15:0] lut_664_table = 16'b1100110011111111;
    wire [3:0] lut_664_select = {
                             in_data[657],
                             in_data[697],
                             in_data[317],
                             in_data[64]};
    
    wire lut_664_out = lut_664_table[lut_664_select];
    
    generate
    if ( USE_REG ) begin : ff_664
        reg   lut_664_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_664_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_664_ff <= lut_664_out;
            end
        end
        
        assign out_data[664] = lut_664_ff;
    end
    else begin : no_ff_664
        assign out_data[664] = lut_664_out;
    end
    endgenerate
    
    
    
    // LUT : 665
    wire [15:0] lut_665_table = 16'b1101010101110001;
    wire [3:0] lut_665_select = {
                             in_data[621],
                             in_data[559],
                             in_data[431],
                             in_data[164]};
    
    wire lut_665_out = lut_665_table[lut_665_select];
    
    generate
    if ( USE_REG ) begin : ff_665
        reg   lut_665_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_665_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_665_ff <= lut_665_out;
            end
        end
        
        assign out_data[665] = lut_665_ff;
    end
    else begin : no_ff_665
        assign out_data[665] = lut_665_out;
    end
    endgenerate
    
    
    
    // LUT : 666
    wire [15:0] lut_666_table = 16'b1010101011111110;
    wire [3:0] lut_666_select = {
                             in_data[41],
                             in_data[771],
                             in_data[243],
                             in_data[116]};
    
    wire lut_666_out = lut_666_table[lut_666_select];
    
    generate
    if ( USE_REG ) begin : ff_666
        reg   lut_666_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_666_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_666_ff <= lut_666_out;
            end
        end
        
        assign out_data[666] = lut_666_ff;
    end
    else begin : no_ff_666
        assign out_data[666] = lut_666_out;
    end
    endgenerate
    
    
    
    // LUT : 667
    wire [15:0] lut_667_table = 16'b1111111111101110;
    wire [3:0] lut_667_select = {
                             in_data[426],
                             in_data[518],
                             in_data[352],
                             in_data[483]};
    
    wire lut_667_out = lut_667_table[lut_667_select];
    
    generate
    if ( USE_REG ) begin : ff_667
        reg   lut_667_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_667_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_667_ff <= lut_667_out;
            end
        end
        
        assign out_data[667] = lut_667_ff;
    end
    else begin : no_ff_667
        assign out_data[667] = lut_667_out;
    end
    endgenerate
    
    
    
    // LUT : 668
    wire [15:0] lut_668_table = 16'b0000000010101010;
    wire [3:0] lut_668_select = {
                             in_data[370],
                             in_data[394],
                             in_data[760],
                             in_data[324]};
    
    wire lut_668_out = lut_668_table[lut_668_select];
    
    generate
    if ( USE_REG ) begin : ff_668
        reg   lut_668_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_668_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_668_ff <= lut_668_out;
            end
        end
        
        assign out_data[668] = lut_668_ff;
    end
    else begin : no_ff_668
        assign out_data[668] = lut_668_out;
    end
    endgenerate
    
    
    
    // LUT : 669
    wire [15:0] lut_669_table = 16'b1101110111001100;
    wire [3:0] lut_669_select = {
                             in_data[242],
                             in_data[111],
                             in_data[99],
                             in_data[172]};
    
    wire lut_669_out = lut_669_table[lut_669_select];
    
    generate
    if ( USE_REG ) begin : ff_669
        reg   lut_669_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_669_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_669_ff <= lut_669_out;
            end
        end
        
        assign out_data[669] = lut_669_ff;
    end
    else begin : no_ff_669
        assign out_data[669] = lut_669_out;
    end
    endgenerate
    
    
    
    // LUT : 670
    wire [15:0] lut_670_table = 16'b1111101010111010;
    wire [3:0] lut_670_select = {
                             in_data[682],
                             in_data[66],
                             in_data[181],
                             in_data[157]};
    
    wire lut_670_out = lut_670_table[lut_670_select];
    
    generate
    if ( USE_REG ) begin : ff_670
        reg   lut_670_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_670_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_670_ff <= lut_670_out;
            end
        end
        
        assign out_data[670] = lut_670_ff;
    end
    else begin : no_ff_670
        assign out_data[670] = lut_670_out;
    end
    endgenerate
    
    
    
    // LUT : 671
    wire [15:0] lut_671_table = 16'b1100110000010001;
    wire [3:0] lut_671_select = {
                             in_data[454],
                             in_data[275],
                             in_data[375],
                             in_data[373]};
    
    wire lut_671_out = lut_671_table[lut_671_select];
    
    generate
    if ( USE_REG ) begin : ff_671
        reg   lut_671_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_671_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_671_ff <= lut_671_out;
            end
        end
        
        assign out_data[671] = lut_671_ff;
    end
    else begin : no_ff_671
        assign out_data[671] = lut_671_out;
    end
    endgenerate
    
    
    
    // LUT : 672
    wire [15:0] lut_672_table = 16'b1111111111111010;
    wire [3:0] lut_672_select = {
                             in_data[70],
                             in_data[711],
                             in_data[312],
                             in_data[750]};
    
    wire lut_672_out = lut_672_table[lut_672_select];
    
    generate
    if ( USE_REG ) begin : ff_672
        reg   lut_672_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_672_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_672_ff <= lut_672_out;
            end
        end
        
        assign out_data[672] = lut_672_ff;
    end
    else begin : no_ff_672
        assign out_data[672] = lut_672_out;
    end
    endgenerate
    
    
    
    // LUT : 673
    wire [15:0] lut_673_table = 16'b0000010001001101;
    wire [3:0] lut_673_select = {
                             in_data[723],
                             in_data[720],
                             in_data[282],
                             in_data[379]};
    
    wire lut_673_out = lut_673_table[lut_673_select];
    
    generate
    if ( USE_REG ) begin : ff_673
        reg   lut_673_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_673_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_673_ff <= lut_673_out;
            end
        end
        
        assign out_data[673] = lut_673_ff;
    end
    else begin : no_ff_673
        assign out_data[673] = lut_673_out;
    end
    endgenerate
    
    
    
    // LUT : 674
    wire [15:0] lut_674_table = 16'b0000000000000101;
    wire [3:0] lut_674_select = {
                             in_data[550],
                             in_data[594],
                             in_data[15],
                             in_data[443]};
    
    wire lut_674_out = lut_674_table[lut_674_select];
    
    generate
    if ( USE_REG ) begin : ff_674
        reg   lut_674_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_674_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_674_ff <= lut_674_out;
            end
        end
        
        assign out_data[674] = lut_674_ff;
    end
    else begin : no_ff_674
        assign out_data[674] = lut_674_out;
    end
    endgenerate
    
    
    
    // LUT : 675
    wire [15:0] lut_675_table = 16'b1111111011111110;
    wire [3:0] lut_675_select = {
                             in_data[82],
                             in_data[75],
                             in_data[194],
                             in_data[632]};
    
    wire lut_675_out = lut_675_table[lut_675_select];
    
    generate
    if ( USE_REG ) begin : ff_675
        reg   lut_675_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_675_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_675_ff <= lut_675_out;
            end
        end
        
        assign out_data[675] = lut_675_ff;
    end
    else begin : no_ff_675
        assign out_data[675] = lut_675_out;
    end
    endgenerate
    
    
    
    // LUT : 676
    wire [15:0] lut_676_table = 16'b0000000000000011;
    wire [3:0] lut_676_select = {
                             in_data[612],
                             in_data[306],
                             in_data[256],
                             in_data[14]};
    
    wire lut_676_out = lut_676_table[lut_676_select];
    
    generate
    if ( USE_REG ) begin : ff_676
        reg   lut_676_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_676_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_676_ff <= lut_676_out;
            end
        end
        
        assign out_data[676] = lut_676_ff;
    end
    else begin : no_ff_676
        assign out_data[676] = lut_676_out;
    end
    endgenerate
    
    
    
    // LUT : 677
    wire [15:0] lut_677_table = 16'b0001000100000000;
    wire [3:0] lut_677_select = {
                             in_data[432],
                             in_data[279],
                             in_data[277],
                             in_data[721]};
    
    wire lut_677_out = lut_677_table[lut_677_select];
    
    generate
    if ( USE_REG ) begin : ff_677
        reg   lut_677_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_677_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_677_ff <= lut_677_out;
            end
        end
        
        assign out_data[677] = lut_677_ff;
    end
    else begin : no_ff_677
        assign out_data[677] = lut_677_out;
    end
    endgenerate
    
    
    
    // LUT : 678
    wire [15:0] lut_678_table = 16'b0000000000010001;
    wire [3:0] lut_678_select = {
                             in_data[226],
                             in_data[757],
                             in_data[87],
                             in_data[738]};
    
    wire lut_678_out = lut_678_table[lut_678_select];
    
    generate
    if ( USE_REG ) begin : ff_678
        reg   lut_678_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_678_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_678_ff <= lut_678_out;
            end
        end
        
        assign out_data[678] = lut_678_ff;
    end
    else begin : no_ff_678
        assign out_data[678] = lut_678_out;
    end
    endgenerate
    
    
    
    // LUT : 679
    wire [15:0] lut_679_table = 16'b0011010100100000;
    wire [3:0] lut_679_select = {
                             in_data[517],
                             in_data[452],
                             in_data[239],
                             in_data[397]};
    
    wire lut_679_out = lut_679_table[lut_679_select];
    
    generate
    if ( USE_REG ) begin : ff_679
        reg   lut_679_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_679_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_679_ff <= lut_679_out;
            end
        end
        
        assign out_data[679] = lut_679_ff;
    end
    else begin : no_ff_679
        assign out_data[679] = lut_679_out;
    end
    endgenerate
    
    
    
    // LUT : 680
    wire [15:0] lut_680_table = 16'b1111111100010000;
    wire [3:0] lut_680_select = {
                             in_data[322],
                             in_data[266],
                             in_data[302],
                             in_data[106]};
    
    wire lut_680_out = lut_680_table[lut_680_select];
    
    generate
    if ( USE_REG ) begin : ff_680
        reg   lut_680_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_680_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_680_ff <= lut_680_out;
            end
        end
        
        assign out_data[680] = lut_680_ff;
    end
    else begin : no_ff_680
        assign out_data[680] = lut_680_out;
    end
    endgenerate
    
    
    
    // LUT : 681
    wire [15:0] lut_681_table = 16'b1100000011111100;
    wire [3:0] lut_681_select = {
                             in_data[643],
                             in_data[231],
                             in_data[142],
                             in_data[672]};
    
    wire lut_681_out = lut_681_table[lut_681_select];
    
    generate
    if ( USE_REG ) begin : ff_681
        reg   lut_681_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_681_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_681_ff <= lut_681_out;
            end
        end
        
        assign out_data[681] = lut_681_ff;
    end
    else begin : no_ff_681
        assign out_data[681] = lut_681_out;
    end
    endgenerate
    
    
    
    // LUT : 682
    wire [15:0] lut_682_table = 16'b1110111011111110;
    wire [3:0] lut_682_select = {
                             in_data[139],
                             in_data[19],
                             in_data[667],
                             in_data[591]};
    
    wire lut_682_out = lut_682_table[lut_682_select];
    
    generate
    if ( USE_REG ) begin : ff_682
        reg   lut_682_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_682_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_682_ff <= lut_682_out;
            end
        end
        
        assign out_data[682] = lut_682_ff;
    end
    else begin : no_ff_682
        assign out_data[682] = lut_682_out;
    end
    endgenerate
    
    
    
    // LUT : 683
    wire [15:0] lut_683_table = 16'b1111111111111110;
    wire [3:0] lut_683_select = {
                             in_data[390],
                             in_data[665],
                             in_data[93],
                             in_data[165]};
    
    wire lut_683_out = lut_683_table[lut_683_select];
    
    generate
    if ( USE_REG ) begin : ff_683
        reg   lut_683_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_683_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_683_ff <= lut_683_out;
            end
        end
        
        assign out_data[683] = lut_683_ff;
    end
    else begin : no_ff_683
        assign out_data[683] = lut_683_out;
    end
    endgenerate
    
    
    
    // LUT : 684
    wire [15:0] lut_684_table = 16'b0000000011111111;
    wire [3:0] lut_684_select = {
                             in_data[606],
                             in_data[297],
                             in_data[167],
                             in_data[380]};
    
    wire lut_684_out = lut_684_table[lut_684_select];
    
    generate
    if ( USE_REG ) begin : ff_684
        reg   lut_684_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_684_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_684_ff <= lut_684_out;
            end
        end
        
        assign out_data[684] = lut_684_ff;
    end
    else begin : no_ff_684
        assign out_data[684] = lut_684_out;
    end
    endgenerate
    
    
    
    // LUT : 685
    wire [15:0] lut_685_table = 16'b1011111110101111;
    wire [3:0] lut_685_select = {
                             in_data[65],
                             in_data[601],
                             in_data[676],
                             in_data[766]};
    
    wire lut_685_out = lut_685_table[lut_685_select];
    
    generate
    if ( USE_REG ) begin : ff_685
        reg   lut_685_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_685_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_685_ff <= lut_685_out;
            end
        end
        
        assign out_data[685] = lut_685_ff;
    end
    else begin : no_ff_685
        assign out_data[685] = lut_685_out;
    end
    endgenerate
    
    
    
    // LUT : 686
    wire [15:0] lut_686_table = 16'b0001000100010001;
    wire [3:0] lut_686_select = {
                             in_data[668],
                             in_data[673],
                             in_data[693],
                             in_data[259]};
    
    wire lut_686_out = lut_686_table[lut_686_select];
    
    generate
    if ( USE_REG ) begin : ff_686
        reg   lut_686_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_686_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_686_ff <= lut_686_out;
            end
        end
        
        assign out_data[686] = lut_686_ff;
    end
    else begin : no_ff_686
        assign out_data[686] = lut_686_out;
    end
    endgenerate
    
    
    
    // LUT : 687
    wire [15:0] lut_687_table = 16'b0000000000101011;
    wire [3:0] lut_687_select = {
                             in_data[415],
                             in_data[283],
                             in_data[234],
                             in_data[748]};
    
    wire lut_687_out = lut_687_table[lut_687_select];
    
    generate
    if ( USE_REG ) begin : ff_687
        reg   lut_687_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_687_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_687_ff <= lut_687_out;
            end
        end
        
        assign out_data[687] = lut_687_ff;
    end
    else begin : no_ff_687
        assign out_data[687] = lut_687_out;
    end
    endgenerate
    
    
    
    // LUT : 688
    wire [15:0] lut_688_table = 16'b0000001000110010;
    wire [3:0] lut_688_select = {
                             in_data[753],
                             in_data[16],
                             in_data[136],
                             in_data[58]};
    
    wire lut_688_out = lut_688_table[lut_688_select];
    
    generate
    if ( USE_REG ) begin : ff_688
        reg   lut_688_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_688_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_688_ff <= lut_688_out;
            end
        end
        
        assign out_data[688] = lut_688_ff;
    end
    else begin : no_ff_688
        assign out_data[688] = lut_688_out;
    end
    endgenerate
    
    
    
    // LUT : 689
    wire [15:0] lut_689_table = 16'b1110111011111110;
    wire [3:0] lut_689_select = {
                             in_data[522],
                             in_data[639],
                             in_data[593],
                             in_data[540]};
    
    wire lut_689_out = lut_689_table[lut_689_select];
    
    generate
    if ( USE_REG ) begin : ff_689
        reg   lut_689_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_689_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_689_ff <= lut_689_out;
            end
        end
        
        assign out_data[689] = lut_689_ff;
    end
    else begin : no_ff_689
        assign out_data[689] = lut_689_out;
    end
    endgenerate
    
    
    
    // LUT : 690
    wire [15:0] lut_690_table = 16'b1101110011011100;
    wire [3:0] lut_690_select = {
                             in_data[57],
                             in_data[177],
                             in_data[122],
                             in_data[103]};
    
    wire lut_690_out = lut_690_table[lut_690_select];
    
    generate
    if ( USE_REG ) begin : ff_690
        reg   lut_690_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_690_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_690_ff <= lut_690_out;
            end
        end
        
        assign out_data[690] = lut_690_ff;
    end
    else begin : no_ff_690
        assign out_data[690] = lut_690_out;
    end
    endgenerate
    
    
    
    // LUT : 691
    wire [15:0] lut_691_table = 16'b0010111100110000;
    wire [3:0] lut_691_select = {
                             in_data[376],
                             in_data[294],
                             in_data[386],
                             in_data[752]};
    
    wire lut_691_out = lut_691_table[lut_691_select];
    
    generate
    if ( USE_REG ) begin : ff_691
        reg   lut_691_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_691_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_691_ff <= lut_691_out;
            end
        end
        
        assign out_data[691] = lut_691_ff;
    end
    else begin : no_ff_691
        assign out_data[691] = lut_691_out;
    end
    endgenerate
    
    
    
    // LUT : 692
    wire [15:0] lut_692_table = 16'b0101010100000101;
    wire [3:0] lut_692_select = {
                             in_data[384],
                             in_data[250],
                             in_data[1],
                             in_data[541]};
    
    wire lut_692_out = lut_692_table[lut_692_select];
    
    generate
    if ( USE_REG ) begin : ff_692
        reg   lut_692_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_692_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_692_ff <= lut_692_out;
            end
        end
        
        assign out_data[692] = lut_692_ff;
    end
    else begin : no_ff_692
        assign out_data[692] = lut_692_out;
    end
    endgenerate
    
    
    
    // LUT : 693
    wire [15:0] lut_693_table = 16'b1111110000111100;
    wire [3:0] lut_693_select = {
                             in_data[604],
                             in_data[650],
                             in_data[570],
                             in_data[590]};
    
    wire lut_693_out = lut_693_table[lut_693_select];
    
    generate
    if ( USE_REG ) begin : ff_693
        reg   lut_693_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_693_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_693_ff <= lut_693_out;
            end
        end
        
        assign out_data[693] = lut_693_ff;
    end
    else begin : no_ff_693
        assign out_data[693] = lut_693_out;
    end
    endgenerate
    
    
    
    // LUT : 694
    wire [15:0] lut_694_table = 16'b1010101011101110;
    wire [3:0] lut_694_select = {
                             in_data[218],
                             in_data[86],
                             in_data[577],
                             in_data[369]};
    
    wire lut_694_out = lut_694_table[lut_694_select];
    
    generate
    if ( USE_REG ) begin : ff_694
        reg   lut_694_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_694_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_694_ff <= lut_694_out;
            end
        end
        
        assign out_data[694] = lut_694_ff;
    end
    else begin : no_ff_694
        assign out_data[694] = lut_694_out;
    end
    endgenerate
    
    
    
    // LUT : 695
    wire [15:0] lut_695_table = 16'b0000101100001111;
    wire [3:0] lut_695_select = {
                             in_data[377],
                             in_data[433],
                             in_data[537],
                             in_data[6]};
    
    wire lut_695_out = lut_695_table[lut_695_select];
    
    generate
    if ( USE_REG ) begin : ff_695
        reg   lut_695_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_695_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_695_ff <= lut_695_out;
            end
        end
        
        assign out_data[695] = lut_695_ff;
    end
    else begin : no_ff_695
        assign out_data[695] = lut_695_out;
    end
    endgenerate
    
    
    
    // LUT : 696
    wire [15:0] lut_696_table = 16'b1101110111001100;
    wire [3:0] lut_696_select = {
                             in_data[300],
                             in_data[4],
                             in_data[608],
                             in_data[76]};
    
    wire lut_696_out = lut_696_table[lut_696_select];
    
    generate
    if ( USE_REG ) begin : ff_696
        reg   lut_696_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_696_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_696_ff <= lut_696_out;
            end
        end
        
        assign out_data[696] = lut_696_ff;
    end
    else begin : no_ff_696
        assign out_data[696] = lut_696_out;
    end
    endgenerate
    
    
    
    // LUT : 697
    wire [15:0] lut_697_table = 16'b1101001111010111;
    wire [3:0] lut_697_select = {
                             in_data[350],
                             in_data[233],
                             in_data[573],
                             in_data[238]};
    
    wire lut_697_out = lut_697_table[lut_697_select];
    
    generate
    if ( USE_REG ) begin : ff_697
        reg   lut_697_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_697_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_697_ff <= lut_697_out;
            end
        end
        
        assign out_data[697] = lut_697_ff;
    end
    else begin : no_ff_697
        assign out_data[697] = lut_697_out;
    end
    endgenerate
    
    
    
    // LUT : 698
    wire [15:0] lut_698_table = 16'b1101110111011101;
    wire [3:0] lut_698_select = {
                             in_data[774],
                             in_data[339],
                             in_data[121],
                             in_data[402]};
    
    wire lut_698_out = lut_698_table[lut_698_select];
    
    generate
    if ( USE_REG ) begin : ff_698
        reg   lut_698_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_698_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_698_ff <= lut_698_out;
            end
        end
        
        assign out_data[698] = lut_698_ff;
    end
    else begin : no_ff_698
        assign out_data[698] = lut_698_out;
    end
    endgenerate
    
    
    
    // LUT : 699
    wire [15:0] lut_699_table = 16'b1111011100111011;
    wire [3:0] lut_699_select = {
                             in_data[610],
                             in_data[493],
                             in_data[574],
                             in_data[214]};
    
    wire lut_699_out = lut_699_table[lut_699_select];
    
    generate
    if ( USE_REG ) begin : ff_699
        reg   lut_699_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_699_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_699_ff <= lut_699_out;
            end
        end
        
        assign out_data[699] = lut_699_ff;
    end
    else begin : no_ff_699
        assign out_data[699] = lut_699_out;
    end
    endgenerate
    
    
    
    // LUT : 700
    wire [15:0] lut_700_table = 16'b1100111110001111;
    wire [3:0] lut_700_select = {
                             in_data[718],
                             in_data[347],
                             in_data[398],
                             in_data[318]};
    
    wire lut_700_out = lut_700_table[lut_700_select];
    
    generate
    if ( USE_REG ) begin : ff_700
        reg   lut_700_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_700_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_700_ff <= lut_700_out;
            end
        end
        
        assign out_data[700] = lut_700_ff;
    end
    else begin : no_ff_700
        assign out_data[700] = lut_700_out;
    end
    endgenerate
    
    
    
    // LUT : 701
    wire [15:0] lut_701_table = 16'b0101000001010101;
    wire [3:0] lut_701_select = {
                             in_data[436],
                             in_data[138],
                             in_data[32],
                             in_data[469]};
    
    wire lut_701_out = lut_701_table[lut_701_select];
    
    generate
    if ( USE_REG ) begin : ff_701
        reg   lut_701_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_701_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_701_ff <= lut_701_out;
            end
        end
        
        assign out_data[701] = lut_701_ff;
    end
    else begin : no_ff_701
        assign out_data[701] = lut_701_out;
    end
    endgenerate
    
    
    
    // LUT : 702
    wire [15:0] lut_702_table = 16'b1111011111010100;
    wire [3:0] lut_702_select = {
                             in_data[217],
                             in_data[656],
                             in_data[160],
                             in_data[240]};
    
    wire lut_702_out = lut_702_table[lut_702_select];
    
    generate
    if ( USE_REG ) begin : ff_702
        reg   lut_702_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_702_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_702_ff <= lut_702_out;
            end
        end
        
        assign out_data[702] = lut_702_ff;
    end
    else begin : no_ff_702
        assign out_data[702] = lut_702_out;
    end
    endgenerate
    
    
    
    // LUT : 703
    wire [15:0] lut_703_table = 16'b1010101010101010;
    wire [3:0] lut_703_select = {
                             in_data[653],
                             in_data[60],
                             in_data[644],
                             in_data[288]};
    
    wire lut_703_out = lut_703_table[lut_703_select];
    
    generate
    if ( USE_REG ) begin : ff_703
        reg   lut_703_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_703_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_703_ff <= lut_703_out;
            end
        end
        
        assign out_data[703] = lut_703_ff;
    end
    else begin : no_ff_703
        assign out_data[703] = lut_703_out;
    end
    endgenerate
    
    
    
    // LUT : 704
    wire [15:0] lut_704_table = 16'b0000000001000101;
    wire [3:0] lut_704_select = {
                             in_data[642],
                             in_data[89],
                             in_data[338],
                             in_data[646]};
    
    wire lut_704_out = lut_704_table[lut_704_select];
    
    generate
    if ( USE_REG ) begin : ff_704
        reg   lut_704_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_704_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_704_ff <= lut_704_out;
            end
        end
        
        assign out_data[704] = lut_704_ff;
    end
    else begin : no_ff_704
        assign out_data[704] = lut_704_out;
    end
    endgenerate
    
    
    
    // LUT : 705
    wire [15:0] lut_705_table = 16'b0101010101000001;
    wire [3:0] lut_705_select = {
                             in_data[199],
                             in_data[499],
                             in_data[156],
                             in_data[178]};
    
    wire lut_705_out = lut_705_table[lut_705_select];
    
    generate
    if ( USE_REG ) begin : ff_705
        reg   lut_705_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_705_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_705_ff <= lut_705_out;
            end
        end
        
        assign out_data[705] = lut_705_ff;
    end
    else begin : no_ff_705
        assign out_data[705] = lut_705_out;
    end
    endgenerate
    
    
    
    // LUT : 706
    wire [15:0] lut_706_table = 16'b1110001001000000;
    wire [3:0] lut_706_select = {
                             in_data[267],
                             in_data[326],
                             in_data[210],
                             in_data[482]};
    
    wire lut_706_out = lut_706_table[lut_706_select];
    
    generate
    if ( USE_REG ) begin : ff_706
        reg   lut_706_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_706_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_706_ff <= lut_706_out;
            end
        end
        
        assign out_data[706] = lut_706_ff;
    end
    else begin : no_ff_706
        assign out_data[706] = lut_706_out;
    end
    endgenerate
    
    
    
    // LUT : 707
    wire [15:0] lut_707_table = 16'b1100000000000011;
    wire [3:0] lut_707_select = {
                             in_data[572],
                             in_data[255],
                             in_data[605],
                             in_data[365]};
    
    wire lut_707_out = lut_707_table[lut_707_select];
    
    generate
    if ( USE_REG ) begin : ff_707
        reg   lut_707_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_707_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_707_ff <= lut_707_out;
            end
        end
        
        assign out_data[707] = lut_707_ff;
    end
    else begin : no_ff_707
        assign out_data[707] = lut_707_out;
    end
    endgenerate
    
    
    
    // LUT : 708
    wire [15:0] lut_708_table = 16'b1111000011110000;
    wire [3:0] lut_708_select = {
                             in_data[684],
                             in_data[180],
                             in_data[0],
                             in_data[779]};
    
    wire lut_708_out = lut_708_table[lut_708_select];
    
    generate
    if ( USE_REG ) begin : ff_708
        reg   lut_708_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_708_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_708_ff <= lut_708_out;
            end
        end
        
        assign out_data[708] = lut_708_ff;
    end
    else begin : no_ff_708
        assign out_data[708] = lut_708_out;
    end
    endgenerate
    
    
    
    // LUT : 709
    wire [15:0] lut_709_table = 16'b0000101000001111;
    wire [3:0] lut_709_select = {
                             in_data[396],
                             in_data[636],
                             in_data[619],
                             in_data[73]};
    
    wire lut_709_out = lut_709_table[lut_709_select];
    
    generate
    if ( USE_REG ) begin : ff_709
        reg   lut_709_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_709_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_709_ff <= lut_709_out;
            end
        end
        
        assign out_data[709] = lut_709_ff;
    end
    else begin : no_ff_709
        assign out_data[709] = lut_709_out;
    end
    endgenerate
    
    
    
    // LUT : 710
    wire [15:0] lut_710_table = 16'b0000101000001010;
    wire [3:0] lut_710_select = {
                             in_data[198],
                             in_data[158],
                             in_data[342],
                             in_data[546]};
    
    wire lut_710_out = lut_710_table[lut_710_select];
    
    generate
    if ( USE_REG ) begin : ff_710
        reg   lut_710_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_710_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_710_ff <= lut_710_out;
            end
        end
        
        assign out_data[710] = lut_710_ff;
    end
    else begin : no_ff_710
        assign out_data[710] = lut_710_out;
    end
    endgenerate
    
    
    
    // LUT : 711
    wire [15:0] lut_711_table = 16'b0101010100010001;
    wire [3:0] lut_711_select = {
                             in_data[252],
                             in_data[728],
                             in_data[113],
                             in_data[554]};
    
    wire lut_711_out = lut_711_table[lut_711_select];
    
    generate
    if ( USE_REG ) begin : ff_711
        reg   lut_711_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_711_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_711_ff <= lut_711_out;
            end
        end
        
        assign out_data[711] = lut_711_ff;
    end
    else begin : no_ff_711
        assign out_data[711] = lut_711_out;
    end
    endgenerate
    
    
    
    // LUT : 712
    wire [15:0] lut_712_table = 16'b0000000001011111;
    wire [3:0] lut_712_select = {
                             in_data[269],
                             in_data[687],
                             in_data[700],
                             in_data[736]};
    
    wire lut_712_out = lut_712_table[lut_712_select];
    
    generate
    if ( USE_REG ) begin : ff_712
        reg   lut_712_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_712_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_712_ff <= lut_712_out;
            end
        end
        
        assign out_data[712] = lut_712_ff;
    end
    else begin : no_ff_712
        assign out_data[712] = lut_712_out;
    end
    endgenerate
    
    
    
    // LUT : 713
    wire [15:0] lut_713_table = 16'b0000000011110010;
    wire [3:0] lut_713_select = {
                             in_data[399],
                             in_data[353],
                             in_data[133],
                             in_data[389]};
    
    wire lut_713_out = lut_713_table[lut_713_select];
    
    generate
    if ( USE_REG ) begin : ff_713
        reg   lut_713_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_713_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_713_ff <= lut_713_out;
            end
        end
        
        assign out_data[713] = lut_713_ff;
    end
    else begin : no_ff_713
        assign out_data[713] = lut_713_out;
    end
    endgenerate
    
    
    
    // LUT : 714
    wire [15:0] lut_714_table = 16'b1111101111111011;
    wire [3:0] lut_714_select = {
                             in_data[314],
                             in_data[72],
                             in_data[183],
                             in_data[595]};
    
    wire lut_714_out = lut_714_table[lut_714_select];
    
    generate
    if ( USE_REG ) begin : ff_714
        reg   lut_714_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_714_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_714_ff <= lut_714_out;
            end
        end
        
        assign out_data[714] = lut_714_ff;
    end
    else begin : no_ff_714
        assign out_data[714] = lut_714_out;
    end
    endgenerate
    
    
    
    // LUT : 715
    wire [15:0] lut_715_table = 16'b1010101010101011;
    wire [3:0] lut_715_select = {
                             in_data[131],
                             in_data[586],
                             in_data[253],
                             in_data[124]};
    
    wire lut_715_out = lut_715_table[lut_715_select];
    
    generate
    if ( USE_REG ) begin : ff_715
        reg   lut_715_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_715_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_715_ff <= lut_715_out;
            end
        end
        
        assign out_data[715] = lut_715_ff;
    end
    else begin : no_ff_715
        assign out_data[715] = lut_715_out;
    end
    endgenerate
    
    
    
    // LUT : 716
    wire [15:0] lut_716_table = 16'b0001000000010111;
    wire [3:0] lut_716_select = {
                             in_data[295],
                             in_data[203],
                             in_data[366],
                             in_data[298]};
    
    wire lut_716_out = lut_716_table[lut_716_select];
    
    generate
    if ( USE_REG ) begin : ff_716
        reg   lut_716_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_716_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_716_ff <= lut_716_out;
            end
        end
        
        assign out_data[716] = lut_716_ff;
    end
    else begin : no_ff_716
        assign out_data[716] = lut_716_out;
    end
    endgenerate
    
    
    
    // LUT : 717
    wire [15:0] lut_717_table = 16'b1111111111111010;
    wire [3:0] lut_717_select = {
                             in_data[175],
                             in_data[710],
                             in_data[685],
                             in_data[584]};
    
    wire lut_717_out = lut_717_table[lut_717_select];
    
    generate
    if ( USE_REG ) begin : ff_717
        reg   lut_717_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_717_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_717_ff <= lut_717_out;
            end
        end
        
        assign out_data[717] = lut_717_ff;
    end
    else begin : no_ff_717
        assign out_data[717] = lut_717_out;
    end
    endgenerate
    
    
    
    // LUT : 718
    wire [15:0] lut_718_table = 16'b0000010100000101;
    wire [3:0] lut_718_select = {
                             in_data[313],
                             in_data[185],
                             in_data[616],
                             in_data[333]};
    
    wire lut_718_out = lut_718_table[lut_718_select];
    
    generate
    if ( USE_REG ) begin : ff_718
        reg   lut_718_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_718_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_718_ff <= lut_718_out;
            end
        end
        
        assign out_data[718] = lut_718_ff;
    end
    else begin : no_ff_718
        assign out_data[718] = lut_718_out;
    end
    endgenerate
    
    
    
    // LUT : 719
    wire [15:0] lut_719_table = 16'b1111111111111110;
    wire [3:0] lut_719_select = {
                             in_data[649],
                             in_data[442],
                             in_data[78],
                             in_data[129]};
    
    wire lut_719_out = lut_719_table[lut_719_select];
    
    generate
    if ( USE_REG ) begin : ff_719
        reg   lut_719_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_719_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_719_ff <= lut_719_out;
            end
        end
        
        assign out_data[719] = lut_719_ff;
    end
    else begin : no_ff_719
        assign out_data[719] = lut_719_out;
    end
    endgenerate
    
    
    
    // LUT : 720
    wire [15:0] lut_720_table = 16'b0000000000000011;
    wire [3:0] lut_720_select = {
                             in_data[263],
                             in_data[337],
                             in_data[741],
                             in_data[501]};
    
    wire lut_720_out = lut_720_table[lut_720_select];
    
    generate
    if ( USE_REG ) begin : ff_720
        reg   lut_720_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_720_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_720_ff <= lut_720_out;
            end
        end
        
        assign out_data[720] = lut_720_ff;
    end
    else begin : no_ff_720
        assign out_data[720] = lut_720_out;
    end
    endgenerate
    
    
    
    // LUT : 721
    wire [15:0] lut_721_table = 16'b1111111110101010;
    wire [3:0] lut_721_select = {
                             in_data[368],
                             in_data[403],
                             in_data[587],
                             in_data[548]};
    
    wire lut_721_out = lut_721_table[lut_721_select];
    
    generate
    if ( USE_REG ) begin : ff_721
        reg   lut_721_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_721_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_721_ff <= lut_721_out;
            end
        end
        
        assign out_data[721] = lut_721_ff;
    end
    else begin : no_ff_721
        assign out_data[721] = lut_721_out;
    end
    endgenerate
    
    
    
    // LUT : 722
    wire [15:0] lut_722_table = 16'b0110111100001111;
    wire [3:0] lut_722_select = {
                             in_data[490],
                             in_data[323],
                             in_data[552],
                             in_data[410]};
    
    wire lut_722_out = lut_722_table[lut_722_select];
    
    generate
    if ( USE_REG ) begin : ff_722
        reg   lut_722_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_722_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_722_ff <= lut_722_out;
            end
        end
        
        assign out_data[722] = lut_722_ff;
    end
    else begin : no_ff_722
        assign out_data[722] = lut_722_out;
    end
    endgenerate
    
    
    
    // LUT : 723
    wire [15:0] lut_723_table = 16'b0000000000010001;
    wire [3:0] lut_723_select = {
                             in_data[479],
                             in_data[671],
                             in_data[563],
                             in_data[340]};
    
    wire lut_723_out = lut_723_table[lut_723_select];
    
    generate
    if ( USE_REG ) begin : ff_723
        reg   lut_723_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_723_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_723_ff <= lut_723_out;
            end
        end
        
        assign out_data[723] = lut_723_ff;
    end
    else begin : no_ff_723
        assign out_data[723] = lut_723_out;
    end
    endgenerate
    
    
    
    // LUT : 724
    wire [15:0] lut_724_table = 16'b1111111100000000;
    wire [3:0] lut_724_select = {
                             in_data[434],
                             in_data[36],
                             in_data[528],
                             in_data[47]};
    
    wire lut_724_out = lut_724_table[lut_724_select];
    
    generate
    if ( USE_REG ) begin : ff_724
        reg   lut_724_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_724_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_724_ff <= lut_724_out;
            end
        end
        
        assign out_data[724] = lut_724_ff;
    end
    else begin : no_ff_724
        assign out_data[724] = lut_724_out;
    end
    endgenerate
    
    
    
    // LUT : 725
    wire [15:0] lut_725_table = 16'b1100000011111110;
    wire [3:0] lut_725_select = {
                             in_data[772],
                             in_data[423],
                             in_data[747],
                             in_data[110]};
    
    wire lut_725_out = lut_725_table[lut_725_select];
    
    generate
    if ( USE_REG ) begin : ff_725
        reg   lut_725_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_725_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_725_ff <= lut_725_out;
            end
        end
        
        assign out_data[725] = lut_725_ff;
    end
    else begin : no_ff_725
        assign out_data[725] = lut_725_out;
    end
    endgenerate
    
    
    
    // LUT : 726
    wire [15:0] lut_726_table = 16'b0000000011110000;
    wire [3:0] lut_726_select = {
                             in_data[221],
                             in_data[489],
                             in_data[363],
                             in_data[633]};
    
    wire lut_726_out = lut_726_table[lut_726_select];
    
    generate
    if ( USE_REG ) begin : ff_726
        reg   lut_726_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_726_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_726_ff <= lut_726_out;
            end
        end
        
        assign out_data[726] = lut_726_ff;
    end
    else begin : no_ff_726
        assign out_data[726] = lut_726_out;
    end
    endgenerate
    
    
    
    // LUT : 727
    wire [15:0] lut_727_table = 16'b1011001010111011;
    wire [3:0] lut_727_select = {
                             in_data[480],
                             in_data[564],
                             in_data[354],
                             in_data[227]};
    
    wire lut_727_out = lut_727_table[lut_727_select];
    
    generate
    if ( USE_REG ) begin : ff_727
        reg   lut_727_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_727_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_727_ff <= lut_727_out;
            end
        end
        
        assign out_data[727] = lut_727_ff;
    end
    else begin : no_ff_727
        assign out_data[727] = lut_727_out;
    end
    endgenerate
    
    
    
    // LUT : 728
    wire [15:0] lut_728_table = 16'b1111110111111101;
    wire [3:0] lut_728_select = {
                             in_data[30],
                             in_data[201],
                             in_data[715],
                             in_data[514]};
    
    wire lut_728_out = lut_728_table[lut_728_select];
    
    generate
    if ( USE_REG ) begin : ff_728
        reg   lut_728_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_728_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_728_ff <= lut_728_out;
            end
        end
        
        assign out_data[728] = lut_728_ff;
    end
    else begin : no_ff_728
        assign out_data[728] = lut_728_out;
    end
    endgenerate
    
    
    
    // LUT : 729
    wire [15:0] lut_729_table = 16'b0000001100000011;
    wire [3:0] lut_729_select = {
                             in_data[189],
                             in_data[425],
                             in_data[712],
                             in_data[688]};
    
    wire lut_729_out = lut_729_table[lut_729_select];
    
    generate
    if ( USE_REG ) begin : ff_729
        reg   lut_729_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_729_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_729_ff <= lut_729_out;
            end
        end
        
        assign out_data[729] = lut_729_ff;
    end
    else begin : no_ff_729
        assign out_data[729] = lut_729_out;
    end
    endgenerate
    
    
    
    // LUT : 730
    wire [15:0] lut_730_table = 16'b0100111111001110;
    wire [3:0] lut_730_select = {
                             in_data[120],
                             in_data[744],
                             in_data[174],
                             in_data[596]};
    
    wire lut_730_out = lut_730_table[lut_730_select];
    
    generate
    if ( USE_REG ) begin : ff_730
        reg   lut_730_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_730_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_730_ff <= lut_730_out;
            end
        end
        
        assign out_data[730] = lut_730_ff;
    end
    else begin : no_ff_730
        assign out_data[730] = lut_730_out;
    end
    endgenerate
    
    
    
    // LUT : 731
    wire [15:0] lut_731_table = 16'b0000000000000001;
    wire [3:0] lut_731_select = {
                             in_data[387],
                             in_data[413],
                             in_data[545],
                             in_data[304]};
    
    wire lut_731_out = lut_731_table[lut_731_select];
    
    generate
    if ( USE_REG ) begin : ff_731
        reg   lut_731_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_731_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_731_ff <= lut_731_out;
            end
        end
        
        assign out_data[731] = lut_731_ff;
    end
    else begin : no_ff_731
        assign out_data[731] = lut_731_out;
    end
    endgenerate
    
    
    
    // LUT : 732
    wire [15:0] lut_732_table = 16'b1111111100100011;
    wire [3:0] lut_732_select = {
                             in_data[293],
                             in_data[731],
                             in_data[492],
                             in_data[470]};
    
    wire lut_732_out = lut_732_table[lut_732_select];
    
    generate
    if ( USE_REG ) begin : ff_732
        reg   lut_732_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_732_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_732_ff <= lut_732_out;
            end
        end
        
        assign out_data[732] = lut_732_ff;
    end
    else begin : no_ff_732
        assign out_data[732] = lut_732_out;
    end
    endgenerate
    
    
    
    // LUT : 733
    wire [15:0] lut_733_table = 16'b1010101010101111;
    wire [3:0] lut_733_select = {
                             in_data[301],
                             in_data[67],
                             in_data[364],
                             in_data[193]};
    
    wire lut_733_out = lut_733_table[lut_733_select];
    
    generate
    if ( USE_REG ) begin : ff_733
        reg   lut_733_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_733_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_733_ff <= lut_733_out;
            end
        end
        
        assign out_data[733] = lut_733_ff;
    end
    else begin : no_ff_733
        assign out_data[733] = lut_733_out;
    end
    endgenerate
    
    
    
    // LUT : 734
    wire [15:0] lut_734_table = 16'b1101110111001100;
    wire [3:0] lut_734_select = {
                             in_data[130],
                             in_data[230],
                             in_data[382],
                             in_data[262]};
    
    wire lut_734_out = lut_734_table[lut_734_select];
    
    generate
    if ( USE_REG ) begin : ff_734
        reg   lut_734_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_734_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_734_ff <= lut_734_out;
            end
        end
        
        assign out_data[734] = lut_734_ff;
    end
    else begin : no_ff_734
        assign out_data[734] = lut_734_out;
    end
    endgenerate
    
    
    
    // LUT : 735
    wire [15:0] lut_735_table = 16'b0000000010101010;
    wire [3:0] lut_735_select = {
                             in_data[118],
                             in_data[420],
                             in_data[54],
                             in_data[289]};
    
    wire lut_735_out = lut_735_table[lut_735_select];
    
    generate
    if ( USE_REG ) begin : ff_735
        reg   lut_735_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_735_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_735_ff <= lut_735_out;
            end
        end
        
        assign out_data[735] = lut_735_ff;
    end
    else begin : no_ff_735
        assign out_data[735] = lut_735_out;
    end
    endgenerate
    
    
    
    // LUT : 736
    wire [15:0] lut_736_table = 16'b0000010000001100;
    wire [3:0] lut_736_select = {
                             in_data[391],
                             in_data[45],
                             in_data[273],
                             in_data[725]};
    
    wire lut_736_out = lut_736_table[lut_736_select];
    
    generate
    if ( USE_REG ) begin : ff_736
        reg   lut_736_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_736_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_736_ff <= lut_736_out;
            end
        end
        
        assign out_data[736] = lut_736_ff;
    end
    else begin : no_ff_736
        assign out_data[736] = lut_736_out;
    end
    endgenerate
    
    
    
    // LUT : 737
    wire [15:0] lut_737_table = 16'b0100010101000101;
    wire [3:0] lut_737_select = {
                             in_data[730],
                             in_data[488],
                             in_data[719],
                             in_data[395]};
    
    wire lut_737_out = lut_737_table[lut_737_select];
    
    generate
    if ( USE_REG ) begin : ff_737
        reg   lut_737_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_737_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_737_ff <= lut_737_out;
            end
        end
        
        assign out_data[737] = lut_737_ff;
    end
    else begin : no_ff_737
        assign out_data[737] = lut_737_out;
    end
    endgenerate
    
    
    
    // LUT : 738
    wire [15:0] lut_738_table = 16'b0011001100110011;
    wire [3:0] lut_738_select = {
                             in_data[95],
                             in_data[274],
                             in_data[463],
                             in_data[477]};
    
    wire lut_738_out = lut_738_table[lut_738_select];
    
    generate
    if ( USE_REG ) begin : ff_738
        reg   lut_738_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_738_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_738_ff <= lut_738_out;
            end
        end
        
        assign out_data[738] = lut_738_ff;
    end
    else begin : no_ff_738
        assign out_data[738] = lut_738_out;
    end
    endgenerate
    
    
    
    // LUT : 739
    wire [15:0] lut_739_table = 16'b0000000000000001;
    wire [3:0] lut_739_select = {
                             in_data[754],
                             in_data[77],
                             in_data[335],
                             in_data[611]};
    
    wire lut_739_out = lut_739_table[lut_739_select];
    
    generate
    if ( USE_REG ) begin : ff_739
        reg   lut_739_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_739_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_739_ff <= lut_739_out;
            end
        end
        
        assign out_data[739] = lut_739_ff;
    end
    else begin : no_ff_739
        assign out_data[739] = lut_739_out;
    end
    endgenerate
    
    
    
    // LUT : 740
    wire [15:0] lut_740_table = 16'b1111110011011100;
    wire [3:0] lut_740_select = {
                             in_data[683],
                             in_data[299],
                             in_data[331],
                             in_data[145]};
    
    wire lut_740_out = lut_740_table[lut_740_select];
    
    generate
    if ( USE_REG ) begin : ff_740
        reg   lut_740_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_740_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_740_ff <= lut_740_out;
            end
        end
        
        assign out_data[740] = lut_740_ff;
    end
    else begin : no_ff_740
        assign out_data[740] = lut_740_out;
    end
    endgenerate
    
    
    
    // LUT : 741
    wire [15:0] lut_741_table = 16'b0000001000001011;
    wire [3:0] lut_741_select = {
                             in_data[600],
                             in_data[544],
                             in_data[68],
                             in_data[290]};
    
    wire lut_741_out = lut_741_table[lut_741_select];
    
    generate
    if ( USE_REG ) begin : ff_741
        reg   lut_741_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_741_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_741_ff <= lut_741_out;
            end
        end
        
        assign out_data[741] = lut_741_ff;
    end
    else begin : no_ff_741
        assign out_data[741] = lut_741_out;
    end
    endgenerate
    
    
    
    // LUT : 742
    wire [15:0] lut_742_table = 16'b1010101011111111;
    wire [3:0] lut_742_select = {
                             in_data[264],
                             in_data[422],
                             in_data[307],
                             in_data[153]};
    
    wire lut_742_out = lut_742_table[lut_742_select];
    
    generate
    if ( USE_REG ) begin : ff_742
        reg   lut_742_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_742_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_742_ff <= lut_742_out;
            end
        end
        
        assign out_data[742] = lut_742_ff;
    end
    else begin : no_ff_742
        assign out_data[742] = lut_742_out;
    end
    endgenerate
    
    
    
    // LUT : 743
    wire [15:0] lut_743_table = 16'b0000001100000011;
    wire [3:0] lut_743_select = {
                             in_data[615],
                             in_data[225],
                             in_data[438],
                             in_data[9]};
    
    wire lut_743_out = lut_743_table[lut_743_select];
    
    generate
    if ( USE_REG ) begin : ff_743
        reg   lut_743_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_743_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_743_ff <= lut_743_out;
            end
        end
        
        assign out_data[743] = lut_743_ff;
    end
    else begin : no_ff_743
        assign out_data[743] = lut_743_out;
    end
    endgenerate
    
    
    
    // LUT : 744
    wire [15:0] lut_744_table = 16'b1111001111110011;
    wire [3:0] lut_744_select = {
                             in_data[703],
                             in_data[742],
                             in_data[406],
                             in_data[626]};
    
    wire lut_744_out = lut_744_table[lut_744_select];
    
    generate
    if ( USE_REG ) begin : ff_744
        reg   lut_744_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_744_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_744_ff <= lut_744_out;
            end
        end
        
        assign out_data[744] = lut_744_ff;
    end
    else begin : no_ff_744
        assign out_data[744] = lut_744_out;
    end
    endgenerate
    
    
    
    // LUT : 745
    wire [15:0] lut_745_table = 16'b1111000011110000;
    wire [3:0] lut_745_select = {
                             in_data[450],
                             in_data[575],
                             in_data[652],
                             in_data[759]};
    
    wire lut_745_out = lut_745_table[lut_745_select];
    
    generate
    if ( USE_REG ) begin : ff_745
        reg   lut_745_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_745_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_745_ff <= lut_745_out;
            end
        end
        
        assign out_data[745] = lut_745_ff;
    end
    else begin : no_ff_745
        assign out_data[745] = lut_745_out;
    end
    endgenerate
    
    
    
    // LUT : 746
    wire [15:0] lut_746_table = 16'b0011000000000111;
    wire [3:0] lut_746_select = {
                             in_data[526],
                             in_data[236],
                             in_data[361],
                             in_data[171]};
    
    wire lut_746_out = lut_746_table[lut_746_select];
    
    generate
    if ( USE_REG ) begin : ff_746
        reg   lut_746_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_746_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_746_ff <= lut_746_out;
            end
        end
        
        assign out_data[746] = lut_746_ff;
    end
    else begin : no_ff_746
        assign out_data[746] = lut_746_out;
    end
    endgenerate
    
    
    
    // LUT : 747
    wire [15:0] lut_747_table = 16'b1101111101001111;
    wire [3:0] lut_747_select = {
                             in_data[666],
                             in_data[349],
                             in_data[679],
                             in_data[100]};
    
    wire lut_747_out = lut_747_table[lut_747_select];
    
    generate
    if ( USE_REG ) begin : ff_747
        reg   lut_747_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_747_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_747_ff <= lut_747_out;
            end
        end
        
        assign out_data[747] = lut_747_ff;
    end
    else begin : no_ff_747
        assign out_data[747] = lut_747_out;
    end
    endgenerate
    
    
    
    // LUT : 748
    wire [15:0] lut_748_table = 16'b1100000011010000;
    wire [3:0] lut_748_select = {
                             in_data[553],
                             in_data[437],
                             in_data[580],
                             in_data[613]};
    
    wire lut_748_out = lut_748_table[lut_748_select];
    
    generate
    if ( USE_REG ) begin : ff_748
        reg   lut_748_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_748_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_748_ff <= lut_748_out;
            end
        end
        
        assign out_data[748] = lut_748_ff;
    end
    else begin : no_ff_748
        assign out_data[748] = lut_748_out;
    end
    endgenerate
    
    
    
    // LUT : 749
    wire [15:0] lut_749_table = 16'b0000000001010000;
    wire [3:0] lut_749_select = {
                             in_data[582],
                             in_data[464],
                             in_data[702],
                             in_data[660]};
    
    wire lut_749_out = lut_749_table[lut_749_select];
    
    generate
    if ( USE_REG ) begin : ff_749
        reg   lut_749_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_749_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_749_ff <= lut_749_out;
            end
        end
        
        assign out_data[749] = lut_749_ff;
    end
    else begin : no_ff_749
        assign out_data[749] = lut_749_out;
    end
    endgenerate
    
    
    
    // LUT : 750
    wire [15:0] lut_750_table = 16'b1110101111001100;
    wire [3:0] lut_750_select = {
                             in_data[458],
                             in_data[371],
                             in_data[461],
                             in_data[362]};
    
    wire lut_750_out = lut_750_table[lut_750_select];
    
    generate
    if ( USE_REG ) begin : ff_750
        reg   lut_750_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_750_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_750_ff <= lut_750_out;
            end
        end
        
        assign out_data[750] = lut_750_ff;
    end
    else begin : no_ff_750
        assign out_data[750] = lut_750_out;
    end
    endgenerate
    
    
    
    // LUT : 751
    wire [15:0] lut_751_table = 16'b0000000000000101;
    wire [3:0] lut_751_select = {
                             in_data[651],
                             in_data[359],
                             in_data[620],
                             in_data[506]};
    
    wire lut_751_out = lut_751_table[lut_751_select];
    
    generate
    if ( USE_REG ) begin : ff_751
        reg   lut_751_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_751_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_751_ff <= lut_751_out;
            end
        end
        
        assign out_data[751] = lut_751_ff;
    end
    else begin : no_ff_751
        assign out_data[751] = lut_751_out;
    end
    endgenerate
    
    
    
    // LUT : 752
    wire [15:0] lut_752_table = 16'b0000000000110010;
    wire [3:0] lut_752_select = {
                             in_data[622],
                             in_data[292],
                             in_data[551],
                             in_data[170]};
    
    wire lut_752_out = lut_752_table[lut_752_select];
    
    generate
    if ( USE_REG ) begin : ff_752
        reg   lut_752_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_752_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_752_ff <= lut_752_out;
            end
        end
        
        assign out_data[752] = lut_752_ff;
    end
    else begin : no_ff_752
        assign out_data[752] = lut_752_out;
    end
    endgenerate
    
    
    
    // LUT : 753
    wire [15:0] lut_753_table = 16'b1111000011110000;
    wire [3:0] lut_753_select = {
                             in_data[59],
                             in_data[268],
                             in_data[560],
                             in_data[235]};
    
    wire lut_753_out = lut_753_table[lut_753_select];
    
    generate
    if ( USE_REG ) begin : ff_753
        reg   lut_753_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_753_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_753_ff <= lut_753_out;
            end
        end
        
        assign out_data[753] = lut_753_ff;
    end
    else begin : no_ff_753
        assign out_data[753] = lut_753_out;
    end
    endgenerate
    
    
    
    // LUT : 754
    wire [15:0] lut_754_table = 16'b0000000000010001;
    wire [3:0] lut_754_select = {
                             in_data[733],
                             in_data[758],
                             in_data[162],
                             in_data[241]};
    
    wire lut_754_out = lut_754_table[lut_754_select];
    
    generate
    if ( USE_REG ) begin : ff_754
        reg   lut_754_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_754_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_754_ff <= lut_754_out;
            end
        end
        
        assign out_data[754] = lut_754_ff;
    end
    else begin : no_ff_754
        assign out_data[754] = lut_754_out;
    end
    endgenerate
    
    
    
    // LUT : 755
    wire [15:0] lut_755_table = 16'b1111111111110000;
    wire [3:0] lut_755_select = {
                             in_data[467],
                             in_data[675],
                             in_data[83],
                             in_data[21]};
    
    wire lut_755_out = lut_755_table[lut_755_select];
    
    generate
    if ( USE_REG ) begin : ff_755
        reg   lut_755_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_755_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_755_ff <= lut_755_out;
            end
        end
        
        assign out_data[755] = lut_755_ff;
    end
    else begin : no_ff_755
        assign out_data[755] = lut_755_out;
    end
    endgenerate
    
    
    
    // LUT : 756
    wire [15:0] lut_756_table = 16'b1111000011111100;
    wire [3:0] lut_756_select = {
                             in_data[276],
                             in_data[466],
                             in_data[530],
                             in_data[699]};
    
    wire lut_756_out = lut_756_table[lut_756_select];
    
    generate
    if ( USE_REG ) begin : ff_756
        reg   lut_756_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_756_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_756_ff <= lut_756_out;
            end
        end
        
        assign out_data[756] = lut_756_ff;
    end
    else begin : no_ff_756
        assign out_data[756] = lut_756_out;
    end
    endgenerate
    
    
    
    // LUT : 757
    wire [15:0] lut_757_table = 16'b1111111100110000;
    wire [3:0] lut_757_select = {
                             in_data[623],
                             in_data[686],
                             in_data[585],
                             in_data[5]};
    
    wire lut_757_out = lut_757_table[lut_757_select];
    
    generate
    if ( USE_REG ) begin : ff_757
        reg   lut_757_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_757_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_757_ff <= lut_757_out;
            end
        end
        
        assign out_data[757] = lut_757_ff;
    end
    else begin : no_ff_757
        assign out_data[757] = lut_757_out;
    end
    endgenerate
    
    
    
    // LUT : 758
    wire [15:0] lut_758_table = 16'b1100110011111110;
    wire [3:0] lut_758_select = {
                             in_data[732],
                             in_data[763],
                             in_data[523],
                             in_data[20]};
    
    wire lut_758_out = lut_758_table[lut_758_select];
    
    generate
    if ( USE_REG ) begin : ff_758
        reg   lut_758_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_758_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_758_ff <= lut_758_out;
            end
        end
        
        assign out_data[758] = lut_758_ff;
    end
    else begin : no_ff_758
        assign out_data[758] = lut_758_out;
    end
    endgenerate
    
    
    
    // LUT : 759
    wire [15:0] lut_759_table = 16'b1111111101010101;
    wire [3:0] lut_759_select = {
                             in_data[722],
                             in_data[765],
                             in_data[780],
                             in_data[599]};
    
    wire lut_759_out = lut_759_table[lut_759_select];
    
    generate
    if ( USE_REG ) begin : ff_759
        reg   lut_759_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_759_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_759_ff <= lut_759_out;
            end
        end
        
        assign out_data[759] = lut_759_ff;
    end
    else begin : no_ff_759
        assign out_data[759] = lut_759_out;
    end
    endgenerate
    
    
    
    // LUT : 760
    wire [15:0] lut_760_table = 16'b1111110011011101;
    wire [3:0] lut_760_select = {
                             in_data[416],
                             in_data[659],
                             in_data[706],
                             in_data[542]};
    
    wire lut_760_out = lut_760_table[lut_760_select];
    
    generate
    if ( USE_REG ) begin : ff_760
        reg   lut_760_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_760_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_760_ff <= lut_760_out;
            end
        end
        
        assign out_data[760] = lut_760_ff;
    end
    else begin : no_ff_760
        assign out_data[760] = lut_760_out;
    end
    endgenerate
    
    
    
    // LUT : 761
    wire [15:0] lut_761_table = 16'b0001000100010001;
    wire [3:0] lut_761_select = {
                             in_data[140],
                             in_data[141],
                             in_data[536],
                             in_data[581]};
    
    wire lut_761_out = lut_761_table[lut_761_select];
    
    generate
    if ( USE_REG ) begin : ff_761
        reg   lut_761_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_761_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_761_ff <= lut_761_out;
            end
        end
        
        assign out_data[761] = lut_761_ff;
    end
    else begin : no_ff_761
        assign out_data[761] = lut_761_out;
    end
    endgenerate
    
    
    
    // LUT : 762
    wire [15:0] lut_762_table = 16'b1010101000100010;
    wire [3:0] lut_762_select = {
                             in_data[664],
                             in_data[114],
                             in_data[108],
                             in_data[655]};
    
    wire lut_762_out = lut_762_table[lut_762_select];
    
    generate
    if ( USE_REG ) begin : ff_762
        reg   lut_762_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_762_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_762_ff <= lut_762_out;
            end
        end
        
        assign out_data[762] = lut_762_ff;
    end
    else begin : no_ff_762
        assign out_data[762] = lut_762_out;
    end
    endgenerate
    
    
    
    // LUT : 763
    wire [15:0] lut_763_table = 16'b0000000011001111;
    wire [3:0] lut_763_select = {
                             in_data[147],
                             in_data[504],
                             in_data[762],
                             in_data[51]};
    
    wire lut_763_out = lut_763_table[lut_763_select];
    
    generate
    if ( USE_REG ) begin : ff_763
        reg   lut_763_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_763_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_763_ff <= lut_763_out;
            end
        end
        
        assign out_data[763] = lut_763_ff;
    end
    else begin : no_ff_763
        assign out_data[763] = lut_763_out;
    end
    endgenerate
    
    
    
    // LUT : 764
    wire [15:0] lut_764_table = 16'b0000101000101011;
    wire [3:0] lut_764_select = {
                             in_data[88],
                             in_data[510],
                             in_data[196],
                             in_data[447]};
    
    wire lut_764_out = lut_764_table[lut_764_select];
    
    generate
    if ( USE_REG ) begin : ff_764
        reg   lut_764_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_764_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_764_ff <= lut_764_out;
            end
        end
        
        assign out_data[764] = lut_764_ff;
    end
    else begin : no_ff_764
        assign out_data[764] = lut_764_out;
    end
    endgenerate
    
    
    
    // LUT : 765
    wire [15:0] lut_765_table = 16'b1111101100001010;
    wire [3:0] lut_765_select = {
                             in_data[498],
                             in_data[691],
                             in_data[117],
                             in_data[330]};
    
    wire lut_765_out = lut_765_table[lut_765_select];
    
    generate
    if ( USE_REG ) begin : ff_765
        reg   lut_765_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_765_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_765_ff <= lut_765_out;
            end
        end
        
        assign out_data[765] = lut_765_ff;
    end
    else begin : no_ff_765
        assign out_data[765] = lut_765_out;
    end
    endgenerate
    
    
    
    // LUT : 766
    wire [15:0] lut_766_table = 16'b0000000000000101;
    wire [3:0] lut_766_select = {
                             in_data[440],
                             in_data[746],
                             in_data[52],
                             in_data[411]};
    
    wire lut_766_out = lut_766_table[lut_766_select];
    
    generate
    if ( USE_REG ) begin : ff_766
        reg   lut_766_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_766_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_766_ff <= lut_766_out;
            end
        end
        
        assign out_data[766] = lut_766_ff;
    end
    else begin : no_ff_766
        assign out_data[766] = lut_766_out;
    end
    endgenerate
    
    
    
    // LUT : 767
    wire [15:0] lut_767_table = 16'b1100110011001100;
    wire [3:0] lut_767_select = {
                             in_data[26],
                             in_data[143],
                             in_data[516],
                             in_data[159]};
    
    wire lut_767_out = lut_767_table[lut_767_select];
    
    generate
    if ( USE_REG ) begin : ff_767
        reg   lut_767_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_767_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_767_ff <= lut_767_out;
            end
        end
        
        assign out_data[767] = lut_767_ff;
    end
    else begin : no_ff_767
        assign out_data[767] = lut_767_out;
    end
    endgenerate
    
    
    
    // LUT : 768
    wire [15:0] lut_768_table = 16'b0100010000001101;
    wire [3:0] lut_768_select = {
                             in_data[182],
                             in_data[569],
                             in_data[271],
                             in_data[692]};
    
    wire lut_768_out = lut_768_table[lut_768_select];
    
    generate
    if ( USE_REG ) begin : ff_768
        reg   lut_768_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_768_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_768_ff <= lut_768_out;
            end
        end
        
        assign out_data[768] = lut_768_ff;
    end
    else begin : no_ff_768
        assign out_data[768] = lut_768_out;
    end
    endgenerate
    
    
    
    // LUT : 769
    wire [15:0] lut_769_table = 16'b0001001100000000;
    wire [3:0] lut_769_select = {
                             in_data[740],
                             in_data[695],
                             in_data[220],
                             in_data[46]};
    
    wire lut_769_out = lut_769_table[lut_769_select];
    
    generate
    if ( USE_REG ) begin : ff_769
        reg   lut_769_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_769_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_769_ff <= lut_769_out;
            end
        end
        
        assign out_data[769] = lut_769_ff;
    end
    else begin : no_ff_769
        assign out_data[769] = lut_769_out;
    end
    endgenerate
    
    
    
    // LUT : 770
    wire [15:0] lut_770_table = 16'b0111111100000001;
    wire [3:0] lut_770_select = {
                             in_data[648],
                             in_data[502],
                             in_data[472],
                             in_data[31]};
    
    wire lut_770_out = lut_770_table[lut_770_select];
    
    generate
    if ( USE_REG ) begin : ff_770
        reg   lut_770_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_770_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_770_ff <= lut_770_out;
            end
        end
        
        assign out_data[770] = lut_770_ff;
    end
    else begin : no_ff_770
        assign out_data[770] = lut_770_out;
    end
    endgenerate
    
    
    
    // LUT : 771
    wire [15:0] lut_771_table = 16'b0000000001010101;
    wire [3:0] lut_771_select = {
                             in_data[97],
                             in_data[80],
                             in_data[583],
                             in_data[212]};
    
    wire lut_771_out = lut_771_table[lut_771_select];
    
    generate
    if ( USE_REG ) begin : ff_771
        reg   lut_771_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_771_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_771_ff <= lut_771_out;
            end
        end
        
        assign out_data[771] = lut_771_ff;
    end
    else begin : no_ff_771
        assign out_data[771] = lut_771_out;
    end
    endgenerate
    
    
    
    // LUT : 772
    wire [15:0] lut_772_table = 16'b1111001111110011;
    wire [3:0] lut_772_select = {
                             in_data[34],
                             in_data[356],
                             in_data[216],
                             in_data[56]};
    
    wire lut_772_out = lut_772_table[lut_772_select];
    
    generate
    if ( USE_REG ) begin : ff_772
        reg   lut_772_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_772_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_772_ff <= lut_772_out;
            end
        end
        
        assign out_data[772] = lut_772_ff;
    end
    else begin : no_ff_772
        assign out_data[772] = lut_772_out;
    end
    endgenerate
    
    
    
    // LUT : 773
    wire [15:0] lut_773_table = 16'b0000000000000101;
    wire [3:0] lut_773_select = {
                             in_data[310],
                             in_data[647],
                             in_data[224],
                             in_data[401]};
    
    wire lut_773_out = lut_773_table[lut_773_select];
    
    generate
    if ( USE_REG ) begin : ff_773
        reg   lut_773_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_773_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_773_ff <= lut_773_out;
            end
        end
        
        assign out_data[773] = lut_773_ff;
    end
    else begin : no_ff_773
        assign out_data[773] = lut_773_out;
    end
    endgenerate
    
    
    
    // LUT : 774
    wire [15:0] lut_774_table = 16'b1000111011001110;
    wire [3:0] lut_774_select = {
                             in_data[478],
                             in_data[126],
                             in_data[681],
                             in_data[678]};
    
    wire lut_774_out = lut_774_table[lut_774_select];
    
    generate
    if ( USE_REG ) begin : ff_774
        reg   lut_774_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_774_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_774_ff <= lut_774_out;
            end
        end
        
        assign out_data[774] = lut_774_ff;
    end
    else begin : no_ff_774
        assign out_data[774] = lut_774_out;
    end
    endgenerate
    
    
    
    // LUT : 775
    wire [15:0] lut_775_table = 16'b1111001100110001;
    wire [3:0] lut_775_select = {
                             in_data[197],
                             in_data[281],
                             in_data[278],
                             in_data[448]};
    
    wire lut_775_out = lut_775_table[lut_775_select];
    
    generate
    if ( USE_REG ) begin : ff_775
        reg   lut_775_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_775_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_775_ff <= lut_775_out;
            end
        end
        
        assign out_data[775] = lut_775_ff;
    end
    else begin : no_ff_775
        assign out_data[775] = lut_775_out;
    end
    endgenerate
    
    
    
    // LUT : 776
    wire [15:0] lut_776_table = 16'b1111101011111010;
    wire [3:0] lut_776_select = {
                             in_data[105],
                             in_data[487],
                             in_data[50],
                             in_data[107]};
    
    wire lut_776_out = lut_776_table[lut_776_select];
    
    generate
    if ( USE_REG ) begin : ff_776
        reg   lut_776_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_776_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_776_ff <= lut_776_out;
            end
        end
        
        assign out_data[776] = lut_776_ff;
    end
    else begin : no_ff_776
        assign out_data[776] = lut_776_out;
    end
    endgenerate
    
    
    
    // LUT : 777
    wire [15:0] lut_777_table = 16'b1111111100110011;
    wire [3:0] lut_777_select = {
                             in_data[446],
                             in_data[309],
                             in_data[321],
                             in_data[776]};
    
    wire lut_777_out = lut_777_table[lut_777_select];
    
    generate
    if ( USE_REG ) begin : ff_777
        reg   lut_777_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_777_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_777_ff <= lut_777_out;
            end
        end
        
        assign out_data[777] = lut_777_ff;
    end
    else begin : no_ff_777
        assign out_data[777] = lut_777_out;
    end
    endgenerate
    
    
    
    // LUT : 778
    wire [15:0] lut_778_table = 16'b1100111011101111;
    wire [3:0] lut_778_select = {
                             in_data[291],
                             in_data[305],
                             in_data[101],
                             in_data[555]};
    
    wire lut_778_out = lut_778_table[lut_778_select];
    
    generate
    if ( USE_REG ) begin : ff_778
        reg   lut_778_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_778_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_778_ff <= lut_778_out;
            end
        end
        
        assign out_data[778] = lut_778_ff;
    end
    else begin : no_ff_778
        assign out_data[778] = lut_778_out;
    end
    endgenerate
    
    
    
    // LUT : 779
    wire [15:0] lut_779_table = 16'b1110111011101110;
    wire [3:0] lut_779_select = {
                             in_data[112],
                             in_data[476],
                             in_data[701],
                             in_data[33]};
    
    wire lut_779_out = lut_779_table[lut_779_select];
    
    generate
    if ( USE_REG ) begin : ff_779
        reg   lut_779_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_779_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_779_ff <= lut_779_out;
            end
        end
        
        assign out_data[779] = lut_779_ff;
    end
    else begin : no_ff_779
        assign out_data[779] = lut_779_out;
    end
    endgenerate
    
    
    
    // LUT : 780
    wire [15:0] lut_780_table = 16'b1111111111111010;
    wire [3:0] lut_780_select = {
                             in_data[202],
                             in_data[424],
                             in_data[775],
                             in_data[609]};
    
    wire lut_780_out = lut_780_table[lut_780_select];
    
    generate
    if ( USE_REG ) begin : ff_780
        reg   lut_780_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_780_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_780_ff <= lut_780_out;
            end
        end
        
        assign out_data[780] = lut_780_ff;
    end
    else begin : no_ff_780
        assign out_data[780] = lut_780_out;
    end
    endgenerate
    
    
    
    // LUT : 781
    wire [15:0] lut_781_table = 16'b0000000000010001;
    wire [3:0] lut_781_select = {
                             in_data[286],
                             in_data[63],
                             in_data[486],
                             in_data[69]};
    
    wire lut_781_out = lut_781_table[lut_781_select];
    
    generate
    if ( USE_REG ) begin : ff_781
        reg   lut_781_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_781_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_781_ff <= lut_781_out;
            end
        end
        
        assign out_data[781] = lut_781_ff;
    end
    else begin : no_ff_781
        assign out_data[781] = lut_781_out;
    end
    endgenerate
    
    
    
    // LUT : 782
    wire [15:0] lut_782_table = 16'b0001000000010001;
    wire [3:0] lut_782_select = {
                             in_data[137],
                             in_data[257],
                             in_data[149],
                             in_data[135]};
    
    wire lut_782_out = lut_782_table[lut_782_select];
    
    generate
    if ( USE_REG ) begin : ff_782
        reg   lut_782_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_782_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_782_ff <= lut_782_out;
            end
        end
        
        assign out_data[782] = lut_782_ff;
    end
    else begin : no_ff_782
        assign out_data[782] = lut_782_out;
    end
    endgenerate
    
    
    
    // LUT : 783
    wire [15:0] lut_783_table = 16'b0000101000001010;
    wire [3:0] lut_783_select = {
                             in_data[475],
                             in_data[258],
                             in_data[18],
                             in_data[405]};
    
    wire lut_783_out = lut_783_table[lut_783_select];
    
    generate
    if ( USE_REG ) begin : ff_783
        reg   lut_783_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_783_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_783_ff <= lut_783_out;
            end
        end
        
        assign out_data[783] = lut_783_ff;
    end
    else begin : no_ff_783
        assign out_data[783] = lut_783_out;
    end
    endgenerate
    
    
    
    // LUT : 784
    wire [15:0] lut_784_table = 16'b1111010100000000;
    wire [3:0] lut_784_select = {
                             in_data[263],
                             in_data[444],
                             in_data[80],
                             in_data[665]};
    
    wire lut_784_out = lut_784_table[lut_784_select];
    
    generate
    if ( USE_REG ) begin : ff_784
        reg   lut_784_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_784_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_784_ff <= lut_784_out;
            end
        end
        
        assign out_data[784] = lut_784_ff;
    end
    else begin : no_ff_784
        assign out_data[784] = lut_784_out;
    end
    endgenerate
    
    
    
    // LUT : 785
    wire [15:0] lut_785_table = 16'b0000000000000101;
    wire [3:0] lut_785_select = {
                             in_data[589],
                             in_data[364],
                             in_data[85],
                             in_data[368]};
    
    wire lut_785_out = lut_785_table[lut_785_select];
    
    generate
    if ( USE_REG ) begin : ff_785
        reg   lut_785_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_785_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_785_ff <= lut_785_out;
            end
        end
        
        assign out_data[785] = lut_785_ff;
    end
    else begin : no_ff_785
        assign out_data[785] = lut_785_out;
    end
    endgenerate
    
    
    
    // LUT : 786
    wire [15:0] lut_786_table = 16'b0000111100001101;
    wire [3:0] lut_786_select = {
                             in_data[500],
                             in_data[314],
                             in_data[119],
                             in_data[265]};
    
    wire lut_786_out = lut_786_table[lut_786_select];
    
    generate
    if ( USE_REG ) begin : ff_786
        reg   lut_786_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_786_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_786_ff <= lut_786_out;
            end
        end
        
        assign out_data[786] = lut_786_ff;
    end
    else begin : no_ff_786
        assign out_data[786] = lut_786_out;
    end
    endgenerate
    
    
    
    // LUT : 787
    wire [15:0] lut_787_table = 16'b0101010101000101;
    wire [3:0] lut_787_select = {
                             in_data[538],
                             in_data[615],
                             in_data[702],
                             in_data[287]};
    
    wire lut_787_out = lut_787_table[lut_787_select];
    
    generate
    if ( USE_REG ) begin : ff_787
        reg   lut_787_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_787_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_787_ff <= lut_787_out;
            end
        end
        
        assign out_data[787] = lut_787_ff;
    end
    else begin : no_ff_787
        assign out_data[787] = lut_787_out;
    end
    endgenerate
    
    
    
    // LUT : 788
    wire [15:0] lut_788_table = 16'b0000010100000101;
    wire [3:0] lut_788_select = {
                             in_data[143],
                             in_data[596],
                             in_data[1],
                             in_data[215]};
    
    wire lut_788_out = lut_788_table[lut_788_select];
    
    generate
    if ( USE_REG ) begin : ff_788
        reg   lut_788_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_788_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_788_ff <= lut_788_out;
            end
        end
        
        assign out_data[788] = lut_788_ff;
    end
    else begin : no_ff_788
        assign out_data[788] = lut_788_out;
    end
    endgenerate
    
    
    
    // LUT : 789
    wire [15:0] lut_789_table = 16'b0000000000000001;
    wire [3:0] lut_789_select = {
                             in_data[565],
                             in_data[528],
                             in_data[172],
                             in_data[231]};
    
    wire lut_789_out = lut_789_table[lut_789_select];
    
    generate
    if ( USE_REG ) begin : ff_789
        reg   lut_789_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_789_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_789_ff <= lut_789_out;
            end
        end
        
        assign out_data[789] = lut_789_ff;
    end
    else begin : no_ff_789
        assign out_data[789] = lut_789_out;
    end
    endgenerate
    
    
    
    // LUT : 790
    wire [15:0] lut_790_table = 16'b0000000011111110;
    wire [3:0] lut_790_select = {
                             in_data[276],
                             in_data[126],
                             in_data[710],
                             in_data[678]};
    
    wire lut_790_out = lut_790_table[lut_790_select];
    
    generate
    if ( USE_REG ) begin : ff_790
        reg   lut_790_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_790_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_790_ff <= lut_790_out;
            end
        end
        
        assign out_data[790] = lut_790_ff;
    end
    else begin : no_ff_790
        assign out_data[790] = lut_790_out;
    end
    endgenerate
    
    
    
    // LUT : 791
    wire [15:0] lut_791_table = 16'b1100000011101100;
    wire [3:0] lut_791_select = {
                             in_data[585],
                             in_data[161],
                             in_data[345],
                             in_data[167]};
    
    wire lut_791_out = lut_791_table[lut_791_select];
    
    generate
    if ( USE_REG ) begin : ff_791
        reg   lut_791_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_791_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_791_ff <= lut_791_out;
            end
        end
        
        assign out_data[791] = lut_791_ff;
    end
    else begin : no_ff_791
        assign out_data[791] = lut_791_out;
    end
    endgenerate
    
    
    
    // LUT : 792
    wire [15:0] lut_792_table = 16'b1010000011111010;
    wire [3:0] lut_792_select = {
                             in_data[691],
                             in_data[525],
                             in_data[36],
                             in_data[633]};
    
    wire lut_792_out = lut_792_table[lut_792_select];
    
    generate
    if ( USE_REG ) begin : ff_792
        reg   lut_792_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_792_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_792_ff <= lut_792_out;
            end
        end
        
        assign out_data[792] = lut_792_ff;
    end
    else begin : no_ff_792
        assign out_data[792] = lut_792_out;
    end
    endgenerate
    
    
    
    // LUT : 793
    wire [15:0] lut_793_table = 16'b1111111110011111;
    wire [3:0] lut_793_select = {
                             in_data[125],
                             in_data[656],
                             in_data[354],
                             in_data[216]};
    
    wire lut_793_out = lut_793_table[lut_793_select];
    
    generate
    if ( USE_REG ) begin : ff_793
        reg   lut_793_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_793_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_793_ff <= lut_793_out;
            end
        end
        
        assign out_data[793] = lut_793_ff;
    end
    else begin : no_ff_793
        assign out_data[793] = lut_793_out;
    end
    endgenerate
    
    
    
    // LUT : 794
    wire [15:0] lut_794_table = 16'b0000000011111111;
    wire [3:0] lut_794_select = {
                             in_data[242],
                             in_data[129],
                             in_data[19],
                             in_data[758]};
    
    wire lut_794_out = lut_794_table[lut_794_select];
    
    generate
    if ( USE_REG ) begin : ff_794
        reg   lut_794_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_794_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_794_ff <= lut_794_out;
            end
        end
        
        assign out_data[794] = lut_794_ff;
    end
    else begin : no_ff_794
        assign out_data[794] = lut_794_out;
    end
    endgenerate
    
    
    
    // LUT : 795
    wire [15:0] lut_795_table = 16'b1111111101000101;
    wire [3:0] lut_795_select = {
                             in_data[708],
                             in_data[616],
                             in_data[554],
                             in_data[372]};
    
    wire lut_795_out = lut_795_table[lut_795_select];
    
    generate
    if ( USE_REG ) begin : ff_795
        reg   lut_795_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_795_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_795_ff <= lut_795_out;
            end
        end
        
        assign out_data[795] = lut_795_ff;
    end
    else begin : no_ff_795
        assign out_data[795] = lut_795_out;
    end
    endgenerate
    
    
    
    // LUT : 796
    wire [15:0] lut_796_table = 16'b0000000000000001;
    wire [3:0] lut_796_select = {
                             in_data[116],
                             in_data[707],
                             in_data[498],
                             in_data[536]};
    
    wire lut_796_out = lut_796_table[lut_796_select];
    
    generate
    if ( USE_REG ) begin : ff_796
        reg   lut_796_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_796_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_796_ff <= lut_796_out;
            end
        end
        
        assign out_data[796] = lut_796_ff;
    end
    else begin : no_ff_796
        assign out_data[796] = lut_796_out;
    end
    endgenerate
    
    
    
    // LUT : 797
    wire [15:0] lut_797_table = 16'b0000000000001100;
    wire [3:0] lut_797_select = {
                             in_data[766],
                             in_data[99],
                             in_data[489],
                             in_data[17]};
    
    wire lut_797_out = lut_797_table[lut_797_select];
    
    generate
    if ( USE_REG ) begin : ff_797
        reg   lut_797_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_797_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_797_ff <= lut_797_out;
            end
        end
        
        assign out_data[797] = lut_797_ff;
    end
    else begin : no_ff_797
        assign out_data[797] = lut_797_out;
    end
    endgenerate
    
    
    
    // LUT : 798
    wire [15:0] lut_798_table = 16'b0101010100000000;
    wire [3:0] lut_798_select = {
                             in_data[625],
                             in_data[617],
                             in_data[141],
                             in_data[748]};
    
    wire lut_798_out = lut_798_table[lut_798_select];
    
    generate
    if ( USE_REG ) begin : ff_798
        reg   lut_798_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_798_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_798_ff <= lut_798_out;
            end
        end
        
        assign out_data[798] = lut_798_ff;
    end
    else begin : no_ff_798
        assign out_data[798] = lut_798_out;
    end
    endgenerate
    
    
    
    // LUT : 799
    wire [15:0] lut_799_table = 16'b0000000000000101;
    wire [3:0] lut_799_select = {
                             in_data[467],
                             in_data[741],
                             in_data[448],
                             in_data[611]};
    
    wire lut_799_out = lut_799_table[lut_799_select];
    
    generate
    if ( USE_REG ) begin : ff_799
        reg   lut_799_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_799_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_799_ff <= lut_799_out;
            end
        end
        
        assign out_data[799] = lut_799_ff;
    end
    else begin : no_ff_799
        assign out_data[799] = lut_799_out;
    end
    endgenerate
    
    
    
    // LUT : 800
    wire [15:0] lut_800_table = 16'b0000000011111111;
    wire [3:0] lut_800_select = {
                             in_data[408],
                             in_data[169],
                             in_data[54],
                             in_data[406]};
    
    wire lut_800_out = lut_800_table[lut_800_select];
    
    generate
    if ( USE_REG ) begin : ff_800
        reg   lut_800_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_800_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_800_ff <= lut_800_out;
            end
        end
        
        assign out_data[800] = lut_800_ff;
    end
    else begin : no_ff_800
        assign out_data[800] = lut_800_out;
    end
    endgenerate
    
    
    
    // LUT : 801
    wire [15:0] lut_801_table = 16'b1100111111001111;
    wire [3:0] lut_801_select = {
                             in_data[251],
                             in_data[155],
                             in_data[356],
                             in_data[739]};
    
    wire lut_801_out = lut_801_table[lut_801_select];
    
    generate
    if ( USE_REG ) begin : ff_801
        reg   lut_801_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_801_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_801_ff <= lut_801_out;
            end
        end
        
        assign out_data[801] = lut_801_ff;
    end
    else begin : no_ff_801
        assign out_data[801] = lut_801_out;
    end
    endgenerate
    
    
    
    // LUT : 802
    wire [15:0] lut_802_table = 16'b0000001100000011;
    wire [3:0] lut_802_select = {
                             in_data[614],
                             in_data[41],
                             in_data[597],
                             in_data[487]};
    
    wire lut_802_out = lut_802_table[lut_802_select];
    
    generate
    if ( USE_REG ) begin : ff_802
        reg   lut_802_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_802_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_802_ff <= lut_802_out;
            end
        end
        
        assign out_data[802] = lut_802_ff;
    end
    else begin : no_ff_802
        assign out_data[802] = lut_802_out;
    end
    endgenerate
    
    
    
    // LUT : 803
    wire [15:0] lut_803_table = 16'b0000000000100011;
    wire [3:0] lut_803_select = {
                             in_data[399],
                             in_data[6],
                             in_data[692],
                             in_data[587]};
    
    wire lut_803_out = lut_803_table[lut_803_select];
    
    generate
    if ( USE_REG ) begin : ff_803
        reg   lut_803_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_803_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_803_ff <= lut_803_out;
            end
        end
        
        assign out_data[803] = lut_803_ff;
    end
    else begin : no_ff_803
        assign out_data[803] = lut_803_out;
    end
    endgenerate
    
    
    
    // LUT : 804
    wire [15:0] lut_804_table = 16'b0000000001000101;
    wire [3:0] lut_804_select = {
                             in_data[325],
                             in_data[299],
                             in_data[51],
                             in_data[501]};
    
    wire lut_804_out = lut_804_table[lut_804_select];
    
    generate
    if ( USE_REG ) begin : ff_804
        reg   lut_804_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_804_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_804_ff <= lut_804_out;
            end
        end
        
        assign out_data[804] = lut_804_ff;
    end
    else begin : no_ff_804
        assign out_data[804] = lut_804_out;
    end
    endgenerate
    
    
    
    // LUT : 805
    wire [15:0] lut_805_table = 16'b0011000011110010;
    wire [3:0] lut_805_select = {
                             in_data[108],
                             in_data[146],
                             in_data[166],
                             in_data[732]};
    
    wire lut_805_out = lut_805_table[lut_805_select];
    
    generate
    if ( USE_REG ) begin : ff_805
        reg   lut_805_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_805_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_805_ff <= lut_805_out;
            end
        end
        
        assign out_data[805] = lut_805_ff;
    end
    else begin : no_ff_805
        assign out_data[805] = lut_805_out;
    end
    endgenerate
    
    
    
    // LUT : 806
    wire [15:0] lut_806_table = 16'b1111111100000000;
    wire [3:0] lut_806_select = {
                             in_data[186],
                             in_data[504],
                             in_data[695],
                             in_data[145]};
    
    wire lut_806_out = lut_806_table[lut_806_select];
    
    generate
    if ( USE_REG ) begin : ff_806
        reg   lut_806_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_806_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_806_ff <= lut_806_out;
            end
        end
        
        assign out_data[806] = lut_806_ff;
    end
    else begin : no_ff_806
        assign out_data[806] = lut_806_out;
    end
    endgenerate
    
    
    
    // LUT : 807
    wire [15:0] lut_807_table = 16'b0000000001000100;
    wire [3:0] lut_807_select = {
                             in_data[734],
                             in_data[420],
                             in_data[603],
                             in_data[738]};
    
    wire lut_807_out = lut_807_table[lut_807_select];
    
    generate
    if ( USE_REG ) begin : ff_807
        reg   lut_807_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_807_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_807_ff <= lut_807_out;
            end
        end
        
        assign out_data[807] = lut_807_ff;
    end
    else begin : no_ff_807
        assign out_data[807] = lut_807_out;
    end
    endgenerate
    
    
    
    // LUT : 808
    wire [15:0] lut_808_table = 16'b1010101010101010;
    wire [3:0] lut_808_select = {
                             in_data[756],
                             in_data[188],
                             in_data[407],
                             in_data[212]};
    
    wire lut_808_out = lut_808_table[lut_808_select];
    
    generate
    if ( USE_REG ) begin : ff_808
        reg   lut_808_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_808_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_808_ff <= lut_808_out;
            end
        end
        
        assign out_data[808] = lut_808_ff;
    end
    else begin : no_ff_808
        assign out_data[808] = lut_808_out;
    end
    endgenerate
    
    
    
    // LUT : 809
    wire [15:0] lut_809_table = 16'b0000000000000001;
    wire [3:0] lut_809_select = {
                             in_data[278],
                             in_data[477],
                             in_data[471],
                             in_data[768]};
    
    wire lut_809_out = lut_809_table[lut_809_select];
    
    generate
    if ( USE_REG ) begin : ff_809
        reg   lut_809_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_809_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_809_ff <= lut_809_out;
            end
        end
        
        assign out_data[809] = lut_809_ff;
    end
    else begin : no_ff_809
        assign out_data[809] = lut_809_out;
    end
    endgenerate
    
    
    
    // LUT : 810
    wire [15:0] lut_810_table = 16'b0011001100110011;
    wire [3:0] lut_810_select = {
                             in_data[105],
                             in_data[754],
                             in_data[295],
                             in_data[514]};
    
    wire lut_810_out = lut_810_table[lut_810_select];
    
    generate
    if ( USE_REG ) begin : ff_810
        reg   lut_810_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_810_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_810_ff <= lut_810_out;
            end
        end
        
        assign out_data[810] = lut_810_ff;
    end
    else begin : no_ff_810
        assign out_data[810] = lut_810_out;
    end
    endgenerate
    
    
    
    // LUT : 811
    wire [15:0] lut_811_table = 16'b0000000011011101;
    wire [3:0] lut_811_select = {
                             in_data[621],
                             in_data[476],
                             in_data[194],
                             in_data[558]};
    
    wire lut_811_out = lut_811_table[lut_811_select];
    
    generate
    if ( USE_REG ) begin : ff_811
        reg   lut_811_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_811_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_811_ff <= lut_811_out;
            end
        end
        
        assign out_data[811] = lut_811_ff;
    end
    else begin : no_ff_811
        assign out_data[811] = lut_811_out;
    end
    endgenerate
    
    
    
    // LUT : 812
    wire [15:0] lut_812_table = 16'b1111111011111110;
    wire [3:0] lut_812_select = {
                             in_data[643],
                             in_data[96],
                             in_data[349],
                             in_data[133]};
    
    wire lut_812_out = lut_812_table[lut_812_select];
    
    generate
    if ( USE_REG ) begin : ff_812
        reg   lut_812_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_812_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_812_ff <= lut_812_out;
            end
        end
        
        assign out_data[812] = lut_812_ff;
    end
    else begin : no_ff_812
        assign out_data[812] = lut_812_out;
    end
    endgenerate
    
    
    
    // LUT : 813
    wire [15:0] lut_813_table = 16'b1000101010111010;
    wire [3:0] lut_813_select = {
                             in_data[666],
                             in_data[256],
                             in_data[348],
                             in_data[327]};
    
    wire lut_813_out = lut_813_table[lut_813_select];
    
    generate
    if ( USE_REG ) begin : ff_813
        reg   lut_813_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_813_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_813_ff <= lut_813_out;
            end
        end
        
        assign out_data[813] = lut_813_ff;
    end
    else begin : no_ff_813
        assign out_data[813] = lut_813_out;
    end
    endgenerate
    
    
    
    // LUT : 814
    wire [15:0] lut_814_table = 16'b1111110111111111;
    wire [3:0] lut_814_select = {
                             in_data[436],
                             in_data[220],
                             in_data[97],
                             in_data[324]};
    
    wire lut_814_out = lut_814_table[lut_814_select];
    
    generate
    if ( USE_REG ) begin : ff_814
        reg   lut_814_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_814_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_814_ff <= lut_814_out;
            end
        end
        
        assign out_data[814] = lut_814_ff;
    end
    else begin : no_ff_814
        assign out_data[814] = lut_814_out;
    end
    endgenerate
    
    
    
    // LUT : 815
    wire [15:0] lut_815_table = 16'b1010101010101110;
    wire [3:0] lut_815_select = {
                             in_data[395],
                             in_data[199],
                             in_data[630],
                             in_data[94]};
    
    wire lut_815_out = lut_815_table[lut_815_select];
    
    generate
    if ( USE_REG ) begin : ff_815
        reg   lut_815_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_815_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_815_ff <= lut_815_out;
            end
        end
        
        assign out_data[815] = lut_815_ff;
    end
    else begin : no_ff_815
        assign out_data[815] = lut_815_out;
    end
    endgenerate
    
    
    
    // LUT : 816
    wire [15:0] lut_816_table = 16'b0011101110101010;
    wire [3:0] lut_816_select = {
                             in_data[268],
                             in_data[660],
                             in_data[534],
                             in_data[456]};
    
    wire lut_816_out = lut_816_table[lut_816_select];
    
    generate
    if ( USE_REG ) begin : ff_816
        reg   lut_816_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_816_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_816_ff <= lut_816_out;
            end
        end
        
        assign out_data[816] = lut_816_ff;
    end
    else begin : no_ff_816
        assign out_data[816] = lut_816_out;
    end
    endgenerate
    
    
    
    // LUT : 817
    wire [15:0] lut_817_table = 16'b0000000011111100;
    wire [3:0] lut_817_select = {
                             in_data[414],
                             in_data[371],
                             in_data[326],
                             in_data[15]};
    
    wire lut_817_out = lut_817_table[lut_817_select];
    
    generate
    if ( USE_REG ) begin : ff_817
        reg   lut_817_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_817_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_817_ff <= lut_817_out;
            end
        end
        
        assign out_data[817] = lut_817_ff;
    end
    else begin : no_ff_817
        assign out_data[817] = lut_817_out;
    end
    endgenerate
    
    
    
    // LUT : 818
    wire [15:0] lut_818_table = 16'b0000111100000101;
    wire [3:0] lut_818_select = {
                             in_data[711],
                             in_data[193],
                             in_data[759],
                             in_data[627]};
    
    wire lut_818_out = lut_818_table[lut_818_select];
    
    generate
    if ( USE_REG ) begin : ff_818
        reg   lut_818_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_818_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_818_ff <= lut_818_out;
            end
        end
        
        assign out_data[818] = lut_818_ff;
    end
    else begin : no_ff_818
        assign out_data[818] = lut_818_out;
    end
    endgenerate
    
    
    
    // LUT : 819
    wire [15:0] lut_819_table = 16'b1111111100010011;
    wire [3:0] lut_819_select = {
                             in_data[446],
                             in_data[168],
                             in_data[382],
                             in_data[699]};
    
    wire lut_819_out = lut_819_table[lut_819_select];
    
    generate
    if ( USE_REG ) begin : ff_819
        reg   lut_819_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_819_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_819_ff <= lut_819_out;
            end
        end
        
        assign out_data[819] = lut_819_ff;
    end
    else begin : no_ff_819
        assign out_data[819] = lut_819_out;
    end
    endgenerate
    
    
    
    // LUT : 820
    wire [15:0] lut_820_table = 16'b0000000000000011;
    wire [3:0] lut_820_select = {
                             in_data[592],
                             in_data[586],
                             in_data[670],
                             in_data[170]};
    
    wire lut_820_out = lut_820_table[lut_820_select];
    
    generate
    if ( USE_REG ) begin : ff_820
        reg   lut_820_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_820_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_820_ff <= lut_820_out;
            end
        end
        
        assign out_data[820] = lut_820_ff;
    end
    else begin : no_ff_820
        assign out_data[820] = lut_820_out;
    end
    endgenerate
    
    
    
    // LUT : 821
    wire [15:0] lut_821_table = 16'b1010101100101011;
    wire [3:0] lut_821_select = {
                             in_data[87],
                             in_data[275],
                             in_data[138],
                             in_data[39]};
    
    wire lut_821_out = lut_821_table[lut_821_select];
    
    generate
    if ( USE_REG ) begin : ff_821
        reg   lut_821_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_821_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_821_ff <= lut_821_out;
            end
        end
        
        assign out_data[821] = lut_821_ff;
    end
    else begin : no_ff_821
        assign out_data[821] = lut_821_out;
    end
    endgenerate
    
    
    
    // LUT : 822
    wire [15:0] lut_822_table = 16'b1111110101000000;
    wire [3:0] lut_822_select = {
                             in_data[239],
                             in_data[594],
                             in_data[679],
                             in_data[78]};
    
    wire lut_822_out = lut_822_table[lut_822_select];
    
    generate
    if ( USE_REG ) begin : ff_822
        reg   lut_822_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_822_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_822_ff <= lut_822_out;
            end
        end
        
        assign out_data[822] = lut_822_ff;
    end
    else begin : no_ff_822
        assign out_data[822] = lut_822_out;
    end
    endgenerate
    
    
    
    // LUT : 823
    wire [15:0] lut_823_table = 16'b0000000000001010;
    wire [3:0] lut_823_select = {
                             in_data[106],
                             in_data[697],
                             in_data[721],
                             in_data[658]};
    
    wire lut_823_out = lut_823_table[lut_823_select];
    
    generate
    if ( USE_REG ) begin : ff_823
        reg   lut_823_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_823_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_823_ff <= lut_823_out;
            end
        end
        
        assign out_data[823] = lut_823_ff;
    end
    else begin : no_ff_823
        assign out_data[823] = lut_823_out;
    end
    endgenerate
    
    
    
    // LUT : 824
    wire [15:0] lut_824_table = 16'b1110111010101010;
    wire [3:0] lut_824_select = {
                             in_data[668],
                             in_data[111],
                             in_data[775],
                             in_data[183]};
    
    wire lut_824_out = lut_824_table[lut_824_select];
    
    generate
    if ( USE_REG ) begin : ff_824
        reg   lut_824_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_824_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_824_ff <= lut_824_out;
            end
        end
        
        assign out_data[824] = lut_824_ff;
    end
    else begin : no_ff_824
        assign out_data[824] = lut_824_out;
    end
    endgenerate
    
    
    
    // LUT : 825
    wire [15:0] lut_825_table = 16'b1000101000101010;
    wire [3:0] lut_825_select = {
                             in_data[75],
                             in_data[472],
                             in_data[132],
                             in_data[655]};
    
    wire lut_825_out = lut_825_table[lut_825_select];
    
    generate
    if ( USE_REG ) begin : ff_825
        reg   lut_825_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_825_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_825_ff <= lut_825_out;
            end
        end
        
        assign out_data[825] = lut_825_ff;
    end
    else begin : no_ff_825
        assign out_data[825] = lut_825_out;
    end
    endgenerate
    
    
    
    // LUT : 826
    wire [15:0] lut_826_table = 16'b1100110011001100;
    wire [3:0] lut_826_select = {
                             in_data[357],
                             in_data[398],
                             in_data[571],
                             in_data[13]};
    
    wire lut_826_out = lut_826_table[lut_826_select];
    
    generate
    if ( USE_REG ) begin : ff_826
        reg   lut_826_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_826_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_826_ff <= lut_826_out;
            end
        end
        
        assign out_data[826] = lut_826_ff;
    end
    else begin : no_ff_826
        assign out_data[826] = lut_826_out;
    end
    endgenerate
    
    
    
    // LUT : 827
    wire [15:0] lut_827_table = 16'b1101111111011101;
    wire [3:0] lut_827_select = {
                             in_data[552],
                             in_data[217],
                             in_data[304],
                             in_data[493]};
    
    wire lut_827_out = lut_827_table[lut_827_select];
    
    generate
    if ( USE_REG ) begin : ff_827
        reg   lut_827_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_827_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_827_ff <= lut_827_out;
            end
        end
        
        assign out_data[827] = lut_827_ff;
    end
    else begin : no_ff_827
        assign out_data[827] = lut_827_out;
    end
    endgenerate
    
    
    
    // LUT : 828
    wire [15:0] lut_828_table = 16'b1101000011110000;
    wire [3:0] lut_828_select = {
                             in_data[67],
                             in_data[431],
                             in_data[599],
                             in_data[203]};
    
    wire lut_828_out = lut_828_table[lut_828_select];
    
    generate
    if ( USE_REG ) begin : ff_828
        reg   lut_828_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_828_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_828_ff <= lut_828_out;
            end
        end
        
        assign out_data[828] = lut_828_ff;
    end
    else begin : no_ff_828
        assign out_data[828] = lut_828_out;
    end
    endgenerate
    
    
    
    // LUT : 829
    wire [15:0] lut_829_table = 16'b0101000000010000;
    wire [3:0] lut_829_select = {
                             in_data[618],
                             in_data[491],
                             in_data[628],
                             in_data[688]};
    
    wire lut_829_out = lut_829_table[lut_829_select];
    
    generate
    if ( USE_REG ) begin : ff_829
        reg   lut_829_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_829_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_829_ff <= lut_829_out;
            end
        end
        
        assign out_data[829] = lut_829_ff;
    end
    else begin : no_ff_829
        assign out_data[829] = lut_829_out;
    end
    endgenerate
    
    
    
    // LUT : 830
    wire [15:0] lut_830_table = 16'b1111001010110000;
    wire [3:0] lut_830_select = {
                             in_data[771],
                             in_data[319],
                             in_data[91],
                             in_data[175]};
    
    wire lut_830_out = lut_830_table[lut_830_select];
    
    generate
    if ( USE_REG ) begin : ff_830
        reg   lut_830_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_830_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_830_ff <= lut_830_out;
            end
        end
        
        assign out_data[830] = lut_830_ff;
    end
    else begin : no_ff_830
        assign out_data[830] = lut_830_out;
    end
    endgenerate
    
    
    
    // LUT : 831
    wire [15:0] lut_831_table = 16'b0000010100000101;
    wire [3:0] lut_831_select = {
                             in_data[689],
                             in_data[257],
                             in_data[765],
                             in_data[274]};
    
    wire lut_831_out = lut_831_table[lut_831_select];
    
    generate
    if ( USE_REG ) begin : ff_831
        reg   lut_831_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_831_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_831_ff <= lut_831_out;
            end
        end
        
        assign out_data[831] = lut_831_ff;
    end
    else begin : no_ff_831
        assign out_data[831] = lut_831_out;
    end
    endgenerate
    
    
    
    // LUT : 832
    wire [15:0] lut_832_table = 16'b0011000100110001;
    wire [3:0] lut_832_select = {
                             in_data[12],
                             in_data[600],
                             in_data[742],
                             in_data[687]};
    
    wire lut_832_out = lut_832_table[lut_832_select];
    
    generate
    if ( USE_REG ) begin : ff_832
        reg   lut_832_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_832_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_832_ff <= lut_832_out;
            end
        end
        
        assign out_data[832] = lut_832_ff;
    end
    else begin : no_ff_832
        assign out_data[832] = lut_832_out;
    end
    endgenerate
    
    
    
    // LUT : 833
    wire [15:0] lut_833_table = 16'b0000111110101110;
    wire [3:0] lut_833_select = {
                             in_data[272],
                             in_data[157],
                             in_data[47],
                             in_data[735]};
    
    wire lut_833_out = lut_833_table[lut_833_select];
    
    generate
    if ( USE_REG ) begin : ff_833
        reg   lut_833_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_833_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_833_ff <= lut_833_out;
            end
        end
        
        assign out_data[833] = lut_833_ff;
    end
    else begin : no_ff_833
        assign out_data[833] = lut_833_out;
    end
    endgenerate
    
    
    
    // LUT : 834
    wire [15:0] lut_834_table = 16'b1110111011111110;
    wire [3:0] lut_834_select = {
                             in_data[777],
                             in_data[550],
                             in_data[177],
                             in_data[123]};
    
    wire lut_834_out = lut_834_table[lut_834_select];
    
    generate
    if ( USE_REG ) begin : ff_834
        reg   lut_834_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_834_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_834_ff <= lut_834_out;
            end
        end
        
        assign out_data[834] = lut_834_ff;
    end
    else begin : no_ff_834
        assign out_data[834] = lut_834_out;
    end
    endgenerate
    
    
    
    // LUT : 835
    wire [15:0] lut_835_table = 16'b0000010000000101;
    wire [3:0] lut_835_select = {
                             in_data[459],
                             in_data[454],
                             in_data[72],
                             in_data[555]};
    
    wire lut_835_out = lut_835_table[lut_835_select];
    
    generate
    if ( USE_REG ) begin : ff_835
        reg   lut_835_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_835_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_835_ff <= lut_835_out;
            end
        end
        
        assign out_data[835] = lut_835_ff;
    end
    else begin : no_ff_835
        assign out_data[835] = lut_835_out;
    end
    endgenerate
    
    
    
    // LUT : 836
    wire [15:0] lut_836_table = 16'b1111001000101011;
    wire [3:0] lut_836_select = {
                             in_data[344],
                             in_data[490],
                             in_data[763],
                             in_data[570]};
    
    wire lut_836_out = lut_836_table[lut_836_select];
    
    generate
    if ( USE_REG ) begin : ff_836
        reg   lut_836_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_836_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_836_ff <= lut_836_out;
            end
        end
        
        assign out_data[836] = lut_836_ff;
    end
    else begin : no_ff_836
        assign out_data[836] = lut_836_out;
    end
    endgenerate
    
    
    
    // LUT : 837
    wire [15:0] lut_837_table = 16'b0101111101011101;
    wire [3:0] lut_837_select = {
                             in_data[416],
                             in_data[680],
                             in_data[542],
                             in_data[264]};
    
    wire lut_837_out = lut_837_table[lut_837_select];
    
    generate
    if ( USE_REG ) begin : ff_837
        reg   lut_837_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_837_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_837_ff <= lut_837_out;
            end
        end
        
        assign out_data[837] = lut_837_ff;
    end
    else begin : no_ff_837
        assign out_data[837] = lut_837_out;
    end
    endgenerate
    
    
    
    // LUT : 838
    wire [15:0] lut_838_table = 16'b0000000011011100;
    wire [3:0] lut_838_select = {
                             in_data[74],
                             in_data[701],
                             in_data[779],
                             in_data[84]};
    
    wire lut_838_out = lut_838_table[lut_838_select];
    
    generate
    if ( USE_REG ) begin : ff_838
        reg   lut_838_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_838_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_838_ff <= lut_838_out;
            end
        end
        
        assign out_data[838] = lut_838_ff;
    end
    else begin : no_ff_838
        assign out_data[838] = lut_838_out;
    end
    endgenerate
    
    
    
    // LUT : 839
    wire [15:0] lut_839_table = 16'b1010101010111011;
    wire [3:0] lut_839_select = {
                             in_data[607],
                             in_data[727],
                             in_data[14],
                             in_data[341]};
    
    wire lut_839_out = lut_839_table[lut_839_select];
    
    generate
    if ( USE_REG ) begin : ff_839
        reg   lut_839_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_839_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_839_ff <= lut_839_out;
            end
        end
        
        assign out_data[839] = lut_839_ff;
    end
    else begin : no_ff_839
        assign out_data[839] = lut_839_out;
    end
    endgenerate
    
    
    
    // LUT : 840
    wire [15:0] lut_840_table = 16'b1111110011111100;
    wire [3:0] lut_840_select = {
                             in_data[417],
                             in_data[153],
                             in_data[44],
                             in_data[73]};
    
    wire lut_840_out = lut_840_table[lut_840_select];
    
    generate
    if ( USE_REG ) begin : ff_840
        reg   lut_840_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_840_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_840_ff <= lut_840_out;
            end
        end
        
        assign out_data[840] = lut_840_ff;
    end
    else begin : no_ff_840
        assign out_data[840] = lut_840_out;
    end
    endgenerate
    
    
    
    // LUT : 841
    wire [15:0] lut_841_table = 16'b0000010100000000;
    wire [3:0] lut_841_select = {
                             in_data[376],
                             in_data[310],
                             in_data[86],
                             in_data[563]};
    
    wire lut_841_out = lut_841_table[lut_841_select];
    
    generate
    if ( USE_REG ) begin : ff_841
        reg   lut_841_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_841_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_841_ff <= lut_841_out;
            end
        end
        
        assign out_data[841] = lut_841_ff;
    end
    else begin : no_ff_841
        assign out_data[841] = lut_841_out;
    end
    endgenerate
    
    
    
    // LUT : 842
    wire [15:0] lut_842_table = 16'b0000000011111111;
    wire [3:0] lut_842_select = {
                             in_data[208],
                             in_data[18],
                             in_data[649],
                             in_data[419]};
    
    wire lut_842_out = lut_842_table[lut_842_select];
    
    generate
    if ( USE_REG ) begin : ff_842
        reg   lut_842_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_842_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_842_ff <= lut_842_out;
            end
        end
        
        assign out_data[842] = lut_842_ff;
    end
    else begin : no_ff_842
        assign out_data[842] = lut_842_out;
    end
    endgenerate
    
    
    
    // LUT : 843
    wire [15:0] lut_843_table = 16'b0000000000110001;
    wire [3:0] lut_843_select = {
                             in_data[45],
                             in_data[88],
                             in_data[450],
                             in_data[158]};
    
    wire lut_843_out = lut_843_table[lut_843_select];
    
    generate
    if ( USE_REG ) begin : ff_843
        reg   lut_843_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_843_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_843_ff <= lut_843_out;
            end
        end
        
        assign out_data[843] = lut_843_ff;
    end
    else begin : no_ff_843
        assign out_data[843] = lut_843_out;
    end
    endgenerate
    
    
    
    // LUT : 844
    wire [15:0] lut_844_table = 16'b0101010101010001;
    wire [3:0] lut_844_select = {
                             in_data[533],
                             in_data[381],
                             in_data[623],
                             in_data[635]};
    
    wire lut_844_out = lut_844_table[lut_844_select];
    
    generate
    if ( USE_REG ) begin : ff_844
        reg   lut_844_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_844_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_844_ff <= lut_844_out;
            end
        end
        
        assign out_data[844] = lut_844_ff;
    end
    else begin : no_ff_844
        assign out_data[844] = lut_844_out;
    end
    endgenerate
    
    
    
    // LUT : 845
    wire [15:0] lut_845_table = 16'b1111111100110011;
    wire [3:0] lut_845_select = {
                             in_data[92],
                             in_data[606],
                             in_data[291],
                             in_data[89]};
    
    wire lut_845_out = lut_845_table[lut_845_select];
    
    generate
    if ( USE_REG ) begin : ff_845
        reg   lut_845_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_845_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_845_ff <= lut_845_out;
            end
        end
        
        assign out_data[845] = lut_845_ff;
    end
    else begin : no_ff_845
        assign out_data[845] = lut_845_out;
    end
    endgenerate
    
    
    
    // LUT : 846
    wire [15:0] lut_846_table = 16'b0100010001000100;
    wire [3:0] lut_846_select = {
                             in_data[21],
                             in_data[253],
                             in_data[405],
                             in_data[537]};
    
    wire lut_846_out = lut_846_table[lut_846_select];
    
    generate
    if ( USE_REG ) begin : ff_846
        reg   lut_846_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_846_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_846_ff <= lut_846_out;
            end
        end
        
        assign out_data[846] = lut_846_ff;
    end
    else begin : no_ff_846
        assign out_data[846] = lut_846_out;
    end
    endgenerate
    
    
    
    // LUT : 847
    wire [15:0] lut_847_table = 16'b0000111100001011;
    wire [3:0] lut_847_select = {
                             in_data[636],
                             in_data[343],
                             in_data[103],
                             in_data[503]};
    
    wire lut_847_out = lut_847_table[lut_847_select];
    
    generate
    if ( USE_REG ) begin : ff_847
        reg   lut_847_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_847_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_847_ff <= lut_847_out;
            end
        end
        
        assign out_data[847] = lut_847_ff;
    end
    else begin : no_ff_847
        assign out_data[847] = lut_847_out;
    end
    endgenerate
    
    
    
    // LUT : 848
    wire [15:0] lut_848_table = 16'b0000000000110011;
    wire [3:0] lut_848_select = {
                             in_data[733],
                             in_data[776],
                             in_data[333],
                             in_data[43]};
    
    wire lut_848_out = lut_848_table[lut_848_select];
    
    generate
    if ( USE_REG ) begin : ff_848
        reg   lut_848_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_848_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_848_ff <= lut_848_out;
            end
        end
        
        assign out_data[848] = lut_848_ff;
    end
    else begin : no_ff_848
        assign out_data[848] = lut_848_out;
    end
    endgenerate
    
    
    
    // LUT : 849
    wire [15:0] lut_849_table = 16'b0000001100000011;
    wire [3:0] lut_849_select = {
                             in_data[79],
                             in_data[207],
                             in_data[64],
                             in_data[57]};
    
    wire lut_849_out = lut_849_table[lut_849_select];
    
    generate
    if ( USE_REG ) begin : ff_849
        reg   lut_849_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_849_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_849_ff <= lut_849_out;
            end
        end
        
        assign out_data[849] = lut_849_ff;
    end
    else begin : no_ff_849
        assign out_data[849] = lut_849_out;
    end
    endgenerate
    
    
    
    // LUT : 850
    wire [15:0] lut_850_table = 16'b0101000011110001;
    wire [3:0] lut_850_select = {
                             in_data[383],
                             in_data[219],
                             in_data[391],
                             in_data[121]};
    
    wire lut_850_out = lut_850_table[lut_850_select];
    
    generate
    if ( USE_REG ) begin : ff_850
        reg   lut_850_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_850_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_850_ff <= lut_850_out;
            end
        end
        
        assign out_data[850] = lut_850_ff;
    end
    else begin : no_ff_850
        assign out_data[850] = lut_850_out;
    end
    endgenerate
    
    
    
    // LUT : 851
    wire [15:0] lut_851_table = 16'b0101010101010101;
    wire [3:0] lut_851_select = {
                             in_data[761],
                             in_data[306],
                             in_data[185],
                             in_data[686]};
    
    wire lut_851_out = lut_851_table[lut_851_select];
    
    generate
    if ( USE_REG ) begin : ff_851
        reg   lut_851_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_851_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_851_ff <= lut_851_out;
            end
        end
        
        assign out_data[851] = lut_851_ff;
    end
    else begin : no_ff_851
        assign out_data[851] = lut_851_out;
    end
    endgenerate
    
    
    
    // LUT : 852
    wire [15:0] lut_852_table = 16'b0000000100010001;
    wire [3:0] lut_852_select = {
                             in_data[159],
                             in_data[548],
                             in_data[524],
                             in_data[180]};
    
    wire lut_852_out = lut_852_table[lut_852_select];
    
    generate
    if ( USE_REG ) begin : ff_852
        reg   lut_852_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_852_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_852_ff <= lut_852_out;
            end
        end
        
        assign out_data[852] = lut_852_ff;
    end
    else begin : no_ff_852
        assign out_data[852] = lut_852_out;
    end
    endgenerate
    
    
    
    // LUT : 853
    wire [15:0] lut_853_table = 16'b0000000000000101;
    wire [3:0] lut_853_select = {
                             in_data[662],
                             in_data[164],
                             in_data[112],
                             in_data[685]};
    
    wire lut_853_out = lut_853_table[lut_853_select];
    
    generate
    if ( USE_REG ) begin : ff_853
        reg   lut_853_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_853_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_853_ff <= lut_853_out;
            end
        end
        
        assign out_data[853] = lut_853_ff;
    end
    else begin : no_ff_853
        assign out_data[853] = lut_853_out;
    end
    endgenerate
    
    
    
    // LUT : 854
    wire [15:0] lut_854_table = 16'b1111000011110000;
    wire [3:0] lut_854_select = {
                             in_data[61],
                             in_data[321],
                             in_data[729],
                             in_data[566]};
    
    wire lut_854_out = lut_854_table[lut_854_select];
    
    generate
    if ( USE_REG ) begin : ff_854
        reg   lut_854_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_854_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_854_ff <= lut_854_out;
            end
        end
        
        assign out_data[854] = lut_854_ff;
    end
    else begin : no_ff_854
        assign out_data[854] = lut_854_out;
    end
    endgenerate
    
    
    
    // LUT : 855
    wire [15:0] lut_855_table = 16'b0000000000101010;
    wire [3:0] lut_855_select = {
                             in_data[329],
                             in_data[359],
                             in_data[465],
                             in_data[403]};
    
    wire lut_855_out = lut_855_table[lut_855_select];
    
    generate
    if ( USE_REG ) begin : ff_855
        reg   lut_855_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_855_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_855_ff <= lut_855_out;
            end
        end
        
        assign out_data[855] = lut_855_ff;
    end
    else begin : no_ff_855
        assign out_data[855] = lut_855_out;
    end
    endgenerate
    
    
    
    // LUT : 856
    wire [15:0] lut_856_table = 16'b0101010101010101;
    wire [3:0] lut_856_select = {
                             in_data[730],
                             in_data[458],
                             in_data[588],
                             in_data[181]};
    
    wire lut_856_out = lut_856_table[lut_856_select];
    
    generate
    if ( USE_REG ) begin : ff_856
        reg   lut_856_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_856_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_856_ff <= lut_856_out;
            end
        end
        
        assign out_data[856] = lut_856_ff;
    end
    else begin : no_ff_856
        assign out_data[856] = lut_856_out;
    end
    endgenerate
    
    
    
    // LUT : 857
    wire [15:0] lut_857_table = 16'b0000101110101010;
    wire [3:0] lut_857_select = {
                             in_data[480],
                             in_data[488],
                             in_data[214],
                             in_data[234]};
    
    wire lut_857_out = lut_857_table[lut_857_select];
    
    generate
    if ( USE_REG ) begin : ff_857
        reg   lut_857_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_857_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_857_ff <= lut_857_out;
            end
        end
        
        assign out_data[857] = lut_857_ff;
    end
    else begin : no_ff_857
        assign out_data[857] = lut_857_out;
    end
    endgenerate
    
    
    
    // LUT : 858
    wire [15:0] lut_858_table = 16'b1111000011110010;
    wire [3:0] lut_858_select = {
                             in_data[745],
                             in_data[497],
                             in_data[361],
                             in_data[437]};
    
    wire lut_858_out = lut_858_table[lut_858_select];
    
    generate
    if ( USE_REG ) begin : ff_858
        reg   lut_858_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_858_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_858_ff <= lut_858_out;
            end
        end
        
        assign out_data[858] = lut_858_ff;
    end
    else begin : no_ff_858
        assign out_data[858] = lut_858_out;
    end
    endgenerate
    
    
    
    // LUT : 859
    wire [15:0] lut_859_table = 16'b0011001100110011;
    wire [3:0] lut_859_select = {
                             in_data[109],
                             in_data[508],
                             in_data[346],
                             in_data[726]};
    
    wire lut_859_out = lut_859_table[lut_859_select];
    
    generate
    if ( USE_REG ) begin : ff_859
        reg   lut_859_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_859_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_859_ff <= lut_859_out;
            end
        end
        
        assign out_data[859] = lut_859_ff;
    end
    else begin : no_ff_859
        assign out_data[859] = lut_859_out;
    end
    endgenerate
    
    
    
    // LUT : 860
    wire [15:0] lut_860_table = 16'b1111111110101010;
    wire [3:0] lut_860_select = {
                             in_data[328],
                             in_data[540],
                             in_data[142],
                             in_data[483]};
    
    wire lut_860_out = lut_860_table[lut_860_select];
    
    generate
    if ( USE_REG ) begin : ff_860
        reg   lut_860_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_860_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_860_ff <= lut_860_out;
            end
        end
        
        assign out_data[860] = lut_860_ff;
    end
    else begin : no_ff_860
        assign out_data[860] = lut_860_out;
    end
    endgenerate
    
    
    
    // LUT : 861
    wire [15:0] lut_861_table = 16'b1011101100100011;
    wire [3:0] lut_861_select = {
                             in_data[475],
                             in_data[0],
                             in_data[62],
                             in_data[674]};
    
    wire lut_861_out = lut_861_table[lut_861_select];
    
    generate
    if ( USE_REG ) begin : ff_861
        reg   lut_861_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_861_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_861_ff <= lut_861_out;
            end
        end
        
        assign out_data[861] = lut_861_ff;
    end
    else begin : no_ff_861
        assign out_data[861] = lut_861_out;
    end
    endgenerate
    
    
    
    // LUT : 862
    wire [15:0] lut_862_table = 16'b0011111110101010;
    wire [3:0] lut_862_select = {
                             in_data[718],
                             in_data[683],
                             in_data[24],
                             in_data[492]};
    
    wire lut_862_out = lut_862_table[lut_862_select];
    
    generate
    if ( USE_REG ) begin : ff_862
        reg   lut_862_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_862_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_862_ff <= lut_862_out;
            end
        end
        
        assign out_data[862] = lut_862_ff;
    end
    else begin : no_ff_862
        assign out_data[862] = lut_862_out;
    end
    endgenerate
    
    
    
    // LUT : 863
    wire [15:0] lut_863_table = 16'b1010101011101110;
    wire [3:0] lut_863_select = {
                             in_data[724],
                             in_data[225],
                             in_data[100],
                             in_data[294]};
    
    wire lut_863_out = lut_863_table[lut_863_select];
    
    generate
    if ( USE_REG ) begin : ff_863
        reg   lut_863_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_863_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_863_ff <= lut_863_out;
            end
        end
        
        assign out_data[863] = lut_863_ff;
    end
    else begin : no_ff_863
        assign out_data[863] = lut_863_out;
    end
    endgenerate
    
    
    
    // LUT : 864
    wire [15:0] lut_864_table = 16'b0000000000001111;
    wire [3:0] lut_864_select = {
                             in_data[95],
                             in_data[574],
                             in_data[530],
                             in_data[139]};
    
    wire lut_864_out = lut_864_table[lut_864_select];
    
    generate
    if ( USE_REG ) begin : ff_864
        reg   lut_864_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_864_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_864_ff <= lut_864_out;
            end
        end
        
        assign out_data[864] = lut_864_ff;
    end
    else begin : no_ff_864
        assign out_data[864] = lut_864_out;
    end
    endgenerate
    
    
    
    // LUT : 865
    wire [15:0] lut_865_table = 16'b1111111110101010;
    wire [3:0] lut_865_select = {
                             in_data[149],
                             in_data[352],
                             in_data[682],
                             in_data[206]};
    
    wire lut_865_out = lut_865_table[lut_865_select];
    
    generate
    if ( USE_REG ) begin : ff_865
        reg   lut_865_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_865_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_865_ff <= lut_865_out;
            end
        end
        
        assign out_data[865] = lut_865_ff;
    end
    else begin : no_ff_865
        assign out_data[865] = lut_865_out;
    end
    endgenerate
    
    
    
    // LUT : 866
    wire [15:0] lut_866_table = 16'b1011111100110011;
    wire [3:0] lut_866_select = {
                             in_data[582],
                             in_data[714],
                             in_data[350],
                             in_data[544]};
    
    wire lut_866_out = lut_866_table[lut_866_select];
    
    generate
    if ( USE_REG ) begin : ff_866
        reg   lut_866_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_866_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_866_ff <= lut_866_out;
            end
        end
        
        assign out_data[866] = lut_866_ff;
    end
    else begin : no_ff_866
        assign out_data[866] = lut_866_out;
    end
    endgenerate
    
    
    
    // LUT : 867
    wire [15:0] lut_867_table = 16'b1100111110001100;
    wire [3:0] lut_867_select = {
                             in_data[93],
                             in_data[165],
                             in_data[466],
                             in_data[53]};
    
    wire lut_867_out = lut_867_table[lut_867_select];
    
    generate
    if ( USE_REG ) begin : ff_867
        reg   lut_867_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_867_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_867_ff <= lut_867_out;
            end
        end
        
        assign out_data[867] = lut_867_ff;
    end
    else begin : no_ff_867
        assign out_data[867] = lut_867_out;
    end
    endgenerate
    
    
    
    // LUT : 868
    wire [15:0] lut_868_table = 16'b1111110011111100;
    wire [3:0] lut_868_select = {
                             in_data[210],
                             in_data[298],
                             in_data[719],
                             in_data[560]};
    
    wire lut_868_out = lut_868_table[lut_868_select];
    
    generate
    if ( USE_REG ) begin : ff_868
        reg   lut_868_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_868_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_868_ff <= lut_868_out;
            end
        end
        
        assign out_data[868] = lut_868_ff;
    end
    else begin : no_ff_868
        assign out_data[868] = lut_868_out;
    end
    endgenerate
    
    
    
    // LUT : 869
    wire [15:0] lut_869_table = 16'b1111101011111010;
    wire [3:0] lut_869_select = {
                             in_data[728],
                             in_data[150],
                             in_data[336],
                             in_data[156]};
    
    wire lut_869_out = lut_869_table[lut_869_select];
    
    generate
    if ( USE_REG ) begin : ff_869
        reg   lut_869_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_869_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_869_ff <= lut_869_out;
            end
        end
        
        assign out_data[869] = lut_869_ff;
    end
    else begin : no_ff_869
        assign out_data[869] = lut_869_out;
    end
    endgenerate
    
    
    
    // LUT : 870
    wire [15:0] lut_870_table = 16'b1010101010101010;
    wire [3:0] lut_870_select = {
                             in_data[66],
                             in_data[81],
                             in_data[33],
                             in_data[315]};
    
    wire lut_870_out = lut_870_table[lut_870_select];
    
    generate
    if ( USE_REG ) begin : ff_870
        reg   lut_870_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_870_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_870_ff <= lut_870_out;
            end
        end
        
        assign out_data[870] = lut_870_ff;
    end
    else begin : no_ff_870
        assign out_data[870] = lut_870_out;
    end
    endgenerate
    
    
    
    // LUT : 871
    wire [15:0] lut_871_table = 16'b0000000100000001;
    wire [3:0] lut_871_select = {
                             in_data[334],
                             in_data[496],
                             in_data[70],
                             in_data[455]};
    
    wire lut_871_out = lut_871_table[lut_871_select];
    
    generate
    if ( USE_REG ) begin : ff_871
        reg   lut_871_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_871_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_871_ff <= lut_871_out;
            end
        end
        
        assign out_data[871] = lut_871_ff;
    end
    else begin : no_ff_871
        assign out_data[871] = lut_871_out;
    end
    endgenerate
    
    
    
    // LUT : 872
    wire [15:0] lut_872_table = 16'b1111000111110001;
    wire [3:0] lut_872_select = {
                             in_data[781],
                             in_data[342],
                             in_data[583],
                             in_data[462]};
    
    wire lut_872_out = lut_872_table[lut_872_select];
    
    generate
    if ( USE_REG ) begin : ff_872
        reg   lut_872_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_872_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_872_ff <= lut_872_out;
            end
        end
        
        assign out_data[872] = lut_872_ff;
    end
    else begin : no_ff_872
        assign out_data[872] = lut_872_out;
    end
    endgenerate
    
    
    
    // LUT : 873
    wire [15:0] lut_873_table = 16'b1111111111111011;
    wire [3:0] lut_873_select = {
                             in_data[284],
                             in_data[178],
                             in_data[572],
                             in_data[740]};
    
    wire lut_873_out = lut_873_table[lut_873_select];
    
    generate
    if ( USE_REG ) begin : ff_873
        reg   lut_873_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_873_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_873_ff <= lut_873_out;
            end
        end
        
        assign out_data[873] = lut_873_ff;
    end
    else begin : no_ff_873
        assign out_data[873] = lut_873_out;
    end
    endgenerate
    
    
    
    // LUT : 874
    wire [15:0] lut_874_table = 16'b1111111100110011;
    wire [3:0] lut_874_select = {
                             in_data[705],
                             in_data[672],
                             in_data[545],
                             in_data[40]};
    
    wire lut_874_out = lut_874_table[lut_874_select];
    
    generate
    if ( USE_REG ) begin : ff_874
        reg   lut_874_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_874_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_874_ff <= lut_874_out;
            end
        end
        
        assign out_data[874] = lut_874_ff;
    end
    else begin : no_ff_874
        assign out_data[874] = lut_874_out;
    end
    endgenerate
    
    
    
    // LUT : 875
    wire [15:0] lut_875_table = 16'b1101110101010100;
    wire [3:0] lut_875_select = {
                             in_data[535],
                             in_data[176],
                             in_data[363],
                             in_data[360]};
    
    wire lut_875_out = lut_875_table[lut_875_select];
    
    generate
    if ( USE_REG ) begin : ff_875
        reg   lut_875_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_875_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_875_ff <= lut_875_out;
            end
        end
        
        assign out_data[875] = lut_875_ff;
    end
    else begin : no_ff_875
        assign out_data[875] = lut_875_out;
    end
    endgenerate
    
    
    
    // LUT : 876
    wire [15:0] lut_876_table = 16'b0101010100000101;
    wire [3:0] lut_876_select = {
                             in_data[227],
                             in_data[522],
                             in_data[657],
                             in_data[204]};
    
    wire lut_876_out = lut_876_table[lut_876_select];
    
    generate
    if ( USE_REG ) begin : ff_876
        reg   lut_876_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_876_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_876_ff <= lut_876_out;
            end
        end
        
        assign out_data[876] = lut_876_ff;
    end
    else begin : no_ff_876
        assign out_data[876] = lut_876_out;
    end
    endgenerate
    
    
    
    // LUT : 877
    wire [15:0] lut_877_table = 16'b1111111011111110;
    wire [3:0] lut_877_select = {
                             in_data[83],
                             in_data[152],
                             in_data[561],
                             in_data[222]};
    
    wire lut_877_out = lut_877_table[lut_877_select];
    
    generate
    if ( USE_REG ) begin : ff_877
        reg   lut_877_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_877_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_877_ff <= lut_877_out;
            end
        end
        
        assign out_data[877] = lut_877_ff;
    end
    else begin : no_ff_877
        assign out_data[877] = lut_877_out;
    end
    endgenerate
    
    
    
    // LUT : 878
    wire [15:0] lut_878_table = 16'b0000010100000101;
    wire [3:0] lut_878_select = {
                             in_data[331],
                             in_data[526],
                             in_data[394],
                             in_data[609]};
    
    wire lut_878_out = lut_878_table[lut_878_select];
    
    generate
    if ( USE_REG ) begin : ff_878
        reg   lut_878_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_878_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_878_ff <= lut_878_out;
            end
        end
        
        assign out_data[878] = lut_878_ff;
    end
    else begin : no_ff_878
        assign out_data[878] = lut_878_out;
    end
    endgenerate
    
    
    
    // LUT : 879
    wire [15:0] lut_879_table = 16'b0101000011111010;
    wire [3:0] lut_879_select = {
                             in_data[367],
                             in_data[470],
                             in_data[113],
                             in_data[452]};
    
    wire lut_879_out = lut_879_table[lut_879_select];
    
    generate
    if ( USE_REG ) begin : ff_879
        reg   lut_879_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_879_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_879_ff <= lut_879_out;
            end
        end
        
        assign out_data[879] = lut_879_ff;
    end
    else begin : no_ff_879
        assign out_data[879] = lut_879_out;
    end
    endgenerate
    
    
    
    // LUT : 880
    wire [15:0] lut_880_table = 16'b0011000000110000;
    wire [3:0] lut_880_select = {
                             in_data[780],
                             in_data[322],
                             in_data[390],
                             in_data[731]};
    
    wire lut_880_out = lut_880_table[lut_880_select];
    
    generate
    if ( USE_REG ) begin : ff_880
        reg   lut_880_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_880_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_880_ff <= lut_880_out;
            end
        end
        
        assign out_data[880] = lut_880_ff;
    end
    else begin : no_ff_880
        assign out_data[880] = lut_880_out;
    end
    endgenerate
    
    
    
    // LUT : 881
    wire [15:0] lut_881_table = 16'b1111111111001101;
    wire [3:0] lut_881_select = {
                             in_data[137],
                             in_data[30],
                             in_data[474],
                             in_data[532]};
    
    wire lut_881_out = lut_881_table[lut_881_select];
    
    generate
    if ( USE_REG ) begin : ff_881
        reg   lut_881_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_881_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_881_ff <= lut_881_out;
            end
        end
        
        assign out_data[881] = lut_881_ff;
    end
    else begin : no_ff_881
        assign out_data[881] = lut_881_out;
    end
    endgenerate
    
    
    
    // LUT : 882
    wire [15:0] lut_882_table = 16'b0000000011001111;
    wire [3:0] lut_882_select = {
                             in_data[218],
                             in_data[353],
                             in_data[418],
                             in_data[279]};
    
    wire lut_882_out = lut_882_table[lut_882_select];
    
    generate
    if ( USE_REG ) begin : ff_882
        reg   lut_882_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_882_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_882_ff <= lut_882_out;
            end
        end
        
        assign out_data[882] = lut_882_ff;
    end
    else begin : no_ff_882
        assign out_data[882] = lut_882_out;
    end
    endgenerate
    
    
    
    // LUT : 883
    wire [15:0] lut_883_table = 16'b0000011100000111;
    wire [3:0] lut_883_select = {
                             in_data[110],
                             in_data[543],
                             in_data[602],
                             in_data[63]};
    
    wire lut_883_out = lut_883_table[lut_883_select];
    
    generate
    if ( USE_REG ) begin : ff_883
        reg   lut_883_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_883_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_883_ff <= lut_883_out;
            end
        end
        
        assign out_data[883] = lut_883_ff;
    end
    else begin : no_ff_883
        assign out_data[883] = lut_883_out;
    end
    endgenerate
    
    
    
    // LUT : 884
    wire [15:0] lut_884_table = 16'b1010101010101010;
    wire [3:0] lut_884_select = {
                             in_data[673],
                             in_data[114],
                             in_data[422],
                             in_data[513]};
    
    wire lut_884_out = lut_884_table[lut_884_select];
    
    generate
    if ( USE_REG ) begin : ff_884
        reg   lut_884_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_884_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_884_ff <= lut_884_out;
            end
        end
        
        assign out_data[884] = lut_884_ff;
    end
    else begin : no_ff_884
        assign out_data[884] = lut_884_out;
    end
    endgenerate
    
    
    
    // LUT : 885
    wire [15:0] lut_885_table = 16'b0000000011101111;
    wire [3:0] lut_885_select = {
                             in_data[486],
                             in_data[261],
                             in_data[440],
                             in_data[421]};
    
    wire lut_885_out = lut_885_table[lut_885_select];
    
    generate
    if ( USE_REG ) begin : ff_885
        reg   lut_885_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_885_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_885_ff <= lut_885_out;
            end
        end
        
        assign out_data[885] = lut_885_ff;
    end
    else begin : no_ff_885
        assign out_data[885] = lut_885_out;
    end
    endgenerate
    
    
    
    // LUT : 886
    wire [15:0] lut_886_table = 16'b0011001100110011;
    wire [3:0] lut_886_select = {
                             in_data[433],
                             in_data[7],
                             in_data[428],
                             in_data[564]};
    
    wire lut_886_out = lut_886_table[lut_886_select];
    
    generate
    if ( USE_REG ) begin : ff_886
        reg   lut_886_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_886_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_886_ff <= lut_886_out;
            end
        end
        
        assign out_data[886] = lut_886_ff;
    end
    else begin : no_ff_886
        assign out_data[886] = lut_886_out;
    end
    endgenerate
    
    
    
    // LUT : 887
    wire [15:0] lut_887_table = 16'b1111111100000000;
    wire [3:0] lut_887_select = {
                             in_data[593],
                             in_data[335],
                             in_data[9],
                             in_data[52]};
    
    wire lut_887_out = lut_887_table[lut_887_select];
    
    generate
    if ( USE_REG ) begin : ff_887
        reg   lut_887_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_887_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_887_ff <= lut_887_out;
            end
        end
        
        assign out_data[887] = lut_887_ff;
    end
    else begin : no_ff_887
        assign out_data[887] = lut_887_out;
    end
    endgenerate
    
    
    
    // LUT : 888
    wire [15:0] lut_888_table = 16'b1111001101110000;
    wire [3:0] lut_888_select = {
                             in_data[610],
                             in_data[460],
                             in_data[259],
                             in_data[478]};
    
    wire lut_888_out = lut_888_table[lut_888_select];
    
    generate
    if ( USE_REG ) begin : ff_888
        reg   lut_888_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_888_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_888_ff <= lut_888_out;
            end
        end
        
        assign out_data[888] = lut_888_ff;
    end
    else begin : no_ff_888
        assign out_data[888] = lut_888_out;
    end
    endgenerate
    
    
    
    // LUT : 889
    wire [15:0] lut_889_table = 16'b1101110111011101;
    wire [3:0] lut_889_select = {
                             in_data[285],
                             in_data[59],
                             in_data[163],
                             in_data[151]};
    
    wire lut_889_out = lut_889_table[lut_889_select];
    
    generate
    if ( USE_REG ) begin : ff_889
        reg   lut_889_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_889_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_889_ff <= lut_889_out;
            end
        end
        
        assign out_data[889] = lut_889_ff;
    end
    else begin : no_ff_889
        assign out_data[889] = lut_889_out;
    end
    endgenerate
    
    
    
    // LUT : 890
    wire [15:0] lut_890_table = 16'b0000000000000101;
    wire [3:0] lut_890_select = {
                             in_data[463],
                             in_data[447],
                             in_data[28],
                             in_data[640]};
    
    wire lut_890_out = lut_890_table[lut_890_select];
    
    generate
    if ( USE_REG ) begin : ff_890
        reg   lut_890_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_890_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_890_ff <= lut_890_out;
            end
        end
        
        assign out_data[890] = lut_890_ff;
    end
    else begin : no_ff_890
        assign out_data[890] = lut_890_out;
    end
    endgenerate
    
    
    
    // LUT : 891
    wire [15:0] lut_891_table = 16'b0100000011011101;
    wire [3:0] lut_891_select = {
                             in_data[388],
                             in_data[307],
                             in_data[42],
                             in_data[198]};
    
    wire lut_891_out = lut_891_table[lut_891_select];
    
    generate
    if ( USE_REG ) begin : ff_891
        reg   lut_891_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_891_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_891_ff <= lut_891_out;
            end
        end
        
        assign out_data[891] = lut_891_ff;
    end
    else begin : no_ff_891
        assign out_data[891] = lut_891_out;
    end
    endgenerate
    
    
    
    // LUT : 892
    wire [15:0] lut_892_table = 16'b1111111110111010;
    wire [3:0] lut_892_select = {
                             in_data[317],
                             in_data[387],
                             in_data[308],
                             in_data[375]};
    
    wire lut_892_out = lut_892_table[lut_892_select];
    
    generate
    if ( USE_REG ) begin : ff_892
        reg   lut_892_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_892_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_892_ff <= lut_892_out;
            end
        end
        
        assign out_data[892] = lut_892_ff;
    end
    else begin : no_ff_892
        assign out_data[892] = lut_892_out;
    end
    endgenerate
    
    
    
    // LUT : 893
    wire [15:0] lut_893_table = 16'b0000101000001111;
    wire [3:0] lut_893_select = {
                             in_data[191],
                             in_data[404],
                             in_data[629],
                             in_data[358]};
    
    wire lut_893_out = lut_893_table[lut_893_select];
    
    generate
    if ( USE_REG ) begin : ff_893
        reg   lut_893_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_893_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_893_ff <= lut_893_out;
            end
        end
        
        assign out_data[893] = lut_893_ff;
    end
    else begin : no_ff_893
        assign out_data[893] = lut_893_out;
    end
    endgenerate
    
    
    
    // LUT : 894
    wire [15:0] lut_894_table = 16'b1100110011001100;
    wire [3:0] lut_894_select = {
                             in_data[26],
                             in_data[144],
                             in_data[634],
                             in_data[288]};
    
    wire lut_894_out = lut_894_table[lut_894_select];
    
    generate
    if ( USE_REG ) begin : ff_894
        reg   lut_894_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_894_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_894_ff <= lut_894_out;
            end
        end
        
        assign out_data[894] = lut_894_ff;
    end
    else begin : no_ff_894
        assign out_data[894] = lut_894_out;
    end
    endgenerate
    
    
    
    // LUT : 895
    wire [15:0] lut_895_table = 16'b1111010111110000;
    wire [3:0] lut_895_select = {
                             in_data[426],
                             in_data[254],
                             in_data[32],
                             in_data[747]};
    
    wire lut_895_out = lut_895_table[lut_895_select];
    
    generate
    if ( USE_REG ) begin : ff_895
        reg   lut_895_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_895_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_895_ff <= lut_895_out;
            end
        end
        
        assign out_data[895] = lut_895_ff;
    end
    else begin : no_ff_895
        assign out_data[895] = lut_895_out;
    end
    endgenerate
    
    
    
    // LUT : 896
    wire [15:0] lut_896_table = 16'b1111111101110000;
    wire [3:0] lut_896_select = {
                             in_data[232],
                             in_data[393],
                             in_data[82],
                             in_data[619]};
    
    wire lut_896_out = lut_896_table[lut_896_select];
    
    generate
    if ( USE_REG ) begin : ff_896
        reg   lut_896_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_896_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_896_ff <= lut_896_out;
            end
        end
        
        assign out_data[896] = lut_896_ff;
    end
    else begin : no_ff_896
        assign out_data[896] = lut_896_out;
    end
    endgenerate
    
    
    
    // LUT : 897
    wire [15:0] lut_897_table = 16'b0111011101100101;
    wire [3:0] lut_897_select = {
                             in_data[485],
                             in_data[620],
                             in_data[102],
                             in_data[270]};
    
    wire lut_897_out = lut_897_table[lut_897_select];
    
    generate
    if ( USE_REG ) begin : ff_897
        reg   lut_897_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_897_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_897_ff <= lut_897_out;
            end
        end
        
        assign out_data[897] = lut_897_ff;
    end
    else begin : no_ff_897
        assign out_data[897] = lut_897_out;
    end
    endgenerate
    
    
    
    // LUT : 898
    wire [15:0] lut_898_table = 16'b0111000111111100;
    wire [3:0] lut_898_select = {
                             in_data[173],
                             in_data[200],
                             in_data[243],
                             in_data[35]};
    
    wire lut_898_out = lut_898_table[lut_898_select];
    
    generate
    if ( USE_REG ) begin : ff_898
        reg   lut_898_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_898_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_898_ff <= lut_898_out;
            end
        end
        
        assign out_data[898] = lut_898_ff;
    end
    else begin : no_ff_898
        assign out_data[898] = lut_898_out;
    end
    endgenerate
    
    
    
    // LUT : 899
    wire [15:0] lut_899_table = 16'b1010000011111111;
    wire [3:0] lut_899_select = {
                             in_data[624],
                             in_data[605],
                             in_data[22],
                             in_data[715]};
    
    wire lut_899_out = lut_899_table[lut_899_select];
    
    generate
    if ( USE_REG ) begin : ff_899
        reg   lut_899_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_899_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_899_ff <= lut_899_out;
            end
        end
        
        assign out_data[899] = lut_899_ff;
    end
    else begin : no_ff_899
        assign out_data[899] = lut_899_out;
    end
    endgenerate
    
    
    
    // LUT : 900
    wire [15:0] lut_900_table = 16'b1111111011101111;
    wire [3:0] lut_900_select = {
                             in_data[397],
                             in_data[575],
                             in_data[622],
                             in_data[709]};
    
    wire lut_900_out = lut_900_table[lut_900_select];
    
    generate
    if ( USE_REG ) begin : ff_900
        reg   lut_900_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_900_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_900_ff <= lut_900_out;
            end
        end
        
        assign out_data[900] = lut_900_ff;
    end
    else begin : no_ff_900
        assign out_data[900] = lut_900_out;
    end
    endgenerate
    
    
    
    // LUT : 901
    wire [15:0] lut_901_table = 16'b1111111111001100;
    wire [3:0] lut_901_select = {
                             in_data[438],
                             in_data[449],
                             in_data[442],
                             in_data[11]};
    
    wire lut_901_out = lut_901_table[lut_901_select];
    
    generate
    if ( USE_REG ) begin : ff_901
        reg   lut_901_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_901_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_901_ff <= lut_901_out;
            end
        end
        
        assign out_data[901] = lut_901_ff;
    end
    else begin : no_ff_901
        assign out_data[901] = lut_901_out;
    end
    endgenerate
    
    
    
    // LUT : 902
    wire [15:0] lut_902_table = 16'b1111111110101010;
    wire [3:0] lut_902_select = {
                             in_data[187],
                             in_data[48],
                             in_data[696],
                             in_data[626]};
    
    wire lut_902_out = lut_902_table[lut_902_select];
    
    generate
    if ( USE_REG ) begin : ff_902
        reg   lut_902_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_902_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_902_ff <= lut_902_out;
            end
        end
        
        assign out_data[902] = lut_902_ff;
    end
    else begin : no_ff_902
        assign out_data[902] = lut_902_out;
    end
    endgenerate
    
    
    
    // LUT : 903
    wire [15:0] lut_903_table = 16'b0000101000001111;
    wire [3:0] lut_903_select = {
                             in_data[774],
                             in_data[521],
                             in_data[65],
                             in_data[230]};
    
    wire lut_903_out = lut_903_table[lut_903_select];
    
    generate
    if ( USE_REG ) begin : ff_903
        reg   lut_903_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_903_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_903_ff <= lut_903_out;
            end
        end
        
        assign out_data[903] = lut_903_ff;
    end
    else begin : no_ff_903
        assign out_data[903] = lut_903_out;
    end
    endgenerate
    
    
    
    // LUT : 904
    wire [15:0] lut_904_table = 16'b1111111111111111;
    wire [3:0] lut_904_select = {
                             in_data[37],
                             in_data[783],
                             in_data[557],
                             in_data[559]};
    
    wire lut_904_out = lut_904_table[lut_904_select];
    
    generate
    if ( USE_REG ) begin : ff_904
        reg   lut_904_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_904_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_904_ff <= lut_904_out;
            end
        end
        
        assign out_data[904] = lut_904_ff;
    end
    else begin : no_ff_904
        assign out_data[904] = lut_904_out;
    end
    endgenerate
    
    
    
    // LUT : 905
    wire [15:0] lut_905_table = 16'b1100111111001100;
    wire [3:0] lut_905_select = {
                             in_data[451],
                             in_data[135],
                             in_data[330],
                             in_data[676]};
    
    wire lut_905_out = lut_905_table[lut_905_select];
    
    generate
    if ( USE_REG ) begin : ff_905
        reg   lut_905_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_905_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_905_ff <= lut_905_out;
            end
        end
        
        assign out_data[905] = lut_905_ff;
    end
    else begin : no_ff_905
        assign out_data[905] = lut_905_out;
    end
    endgenerate
    
    
    
    // LUT : 906
    wire [15:0] lut_906_table = 16'b0101011100000000;
    wire [3:0] lut_906_select = {
                             in_data[303],
                             in_data[195],
                             in_data[197],
                             in_data[772]};
    
    wire lut_906_out = lut_906_table[lut_906_select];
    
    generate
    if ( USE_REG ) begin : ff_906
        reg   lut_906_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_906_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_906_ff <= lut_906_out;
            end
        end
        
        assign out_data[906] = lut_906_ff;
    end
    else begin : no_ff_906
        assign out_data[906] = lut_906_out;
    end
    endgenerate
    
    
    
    // LUT : 907
    wire [15:0] lut_907_table = 16'b1111000011110000;
    wire [3:0] lut_907_select = {
                             in_data[577],
                             in_data[659],
                             in_data[693],
                             in_data[505]};
    
    wire lut_907_out = lut_907_table[lut_907_select];
    
    generate
    if ( USE_REG ) begin : ff_907
        reg   lut_907_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_907_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_907_ff <= lut_907_out;
            end
        end
        
        assign out_data[907] = lut_907_ff;
    end
    else begin : no_ff_907
        assign out_data[907] = lut_907_out;
    end
    endgenerate
    
    
    
    // LUT : 908
    wire [15:0] lut_908_table = 16'b1111111111110000;
    wire [3:0] lut_908_select = {
                             in_data[339],
                             in_data[297],
                             in_data[671],
                             in_data[631]};
    
    wire lut_908_out = lut_908_table[lut_908_select];
    
    generate
    if ( USE_REG ) begin : ff_908
        reg   lut_908_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_908_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_908_ff <= lut_908_out;
            end
        end
        
        assign out_data[908] = lut_908_ff;
    end
    else begin : no_ff_908
        assign out_data[908] = lut_908_out;
    end
    endgenerate
    
    
    
    // LUT : 909
    wire [15:0] lut_909_table = 16'b1111111101110000;
    wire [3:0] lut_909_select = {
                             in_data[743],
                             in_data[240],
                             in_data[647],
                             in_data[373]};
    
    wire lut_909_out = lut_909_table[lut_909_select];
    
    generate
    if ( USE_REG ) begin : ff_909
        reg   lut_909_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_909_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_909_ff <= lut_909_out;
            end
        end
        
        assign out_data[909] = lut_909_ff;
    end
    else begin : no_ff_909
        assign out_data[909] = lut_909_out;
    end
    endgenerate
    
    
    
    // LUT : 910
    wire [15:0] lut_910_table = 16'b1100110011101111;
    wire [3:0] lut_910_select = {
                             in_data[128],
                             in_data[590],
                             in_data[716],
                             in_data[365]};
    
    wire lut_910_out = lut_910_table[lut_910_select];
    
    generate
    if ( USE_REG ) begin : ff_910
        reg   lut_910_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_910_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_910_ff <= lut_910_out;
            end
        end
        
        assign out_data[910] = lut_910_ff;
    end
    else begin : no_ff_910
        assign out_data[910] = lut_910_out;
    end
    endgenerate
    
    
    
    // LUT : 911
    wire [15:0] lut_911_table = 16'b0000000011111111;
    wire [3:0] lut_911_select = {
                             in_data[205],
                             in_data[309],
                             in_data[10],
                             in_data[494]};
    
    wire lut_911_out = lut_911_table[lut_911_select];
    
    generate
    if ( USE_REG ) begin : ff_911
        reg   lut_911_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_911_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_911_ff <= lut_911_out;
            end
        end
        
        assign out_data[911] = lut_911_ff;
    end
    else begin : no_ff_911
        assign out_data[911] = lut_911_out;
    end
    endgenerate
    
    
    
    // LUT : 912
    wire [15:0] lut_912_table = 16'b0000000011110001;
    wire [3:0] lut_912_select = {
                             in_data[104],
                             in_data[512],
                             in_data[652],
                             in_data[591]};
    
    wire lut_912_out = lut_912_table[lut_912_select];
    
    generate
    if ( USE_REG ) begin : ff_912
        reg   lut_912_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_912_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_912_ff <= lut_912_out;
            end
        end
        
        assign out_data[912] = lut_912_ff;
    end
    else begin : no_ff_912
        assign out_data[912] = lut_912_out;
    end
    endgenerate
    
    
    
    // LUT : 913
    wire [15:0] lut_913_table = 16'b0011101100110011;
    wire [3:0] lut_913_select = {
                             in_data[764],
                             in_data[312],
                             in_data[461],
                             in_data[179]};
    
    wire lut_913_out = lut_913_table[lut_913_select];
    
    generate
    if ( USE_REG ) begin : ff_913
        reg   lut_913_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_913_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_913_ff <= lut_913_out;
            end
        end
        
        assign out_data[913] = lut_913_ff;
    end
    else begin : no_ff_913
        assign out_data[913] = lut_913_out;
    end
    endgenerate
    
    
    
    // LUT : 914
    wire [15:0] lut_914_table = 16'b0001000100010001;
    wire [3:0] lut_914_select = {
                             in_data[644],
                             in_data[663],
                             in_data[190],
                             in_data[370]};
    
    wire lut_914_out = lut_914_table[lut_914_select];
    
    generate
    if ( USE_REG ) begin : ff_914
        reg   lut_914_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_914_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_914_ff <= lut_914_out;
            end
        end
        
        assign out_data[914] = lut_914_ff;
    end
    else begin : no_ff_914
        assign out_data[914] = lut_914_out;
    end
    endgenerate
    
    
    
    // LUT : 915
    wire [15:0] lut_915_table = 16'b0000010000001100;
    wire [3:0] lut_915_select = {
                             in_data[384],
                             in_data[651],
                             in_data[271],
                             in_data[736]};
    
    wire lut_915_out = lut_915_table[lut_915_select];
    
    generate
    if ( USE_REG ) begin : ff_915
        reg   lut_915_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_915_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_915_ff <= lut_915_out;
            end
        end
        
        assign out_data[915] = lut_915_ff;
    end
    else begin : no_ff_915
        assign out_data[915] = lut_915_out;
    end
    endgenerate
    
    
    
    // LUT : 916
    wire [15:0] lut_916_table = 16'b0011001000110001;
    wire [3:0] lut_916_select = {
                             in_data[27],
                             in_data[499],
                             in_data[713],
                             in_data[29]};
    
    wire lut_916_out = lut_916_table[lut_916_select];
    
    generate
    if ( USE_REG ) begin : ff_916
        reg   lut_916_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_916_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_916_ff <= lut_916_out;
            end
        end
        
        assign out_data[916] = lut_916_ff;
    end
    else begin : no_ff_916
        assign out_data[916] = lut_916_out;
    end
    endgenerate
    
    
    
    // LUT : 917
    wire [15:0] lut_917_table = 16'b0111001100000011;
    wire [3:0] lut_917_select = {
                             in_data[576],
                             in_data[516],
                             in_data[546],
                             in_data[767]};
    
    wire lut_917_out = lut_917_table[lut_917_select];
    
    generate
    if ( USE_REG ) begin : ff_917
        reg   lut_917_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_917_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_917_ff <= lut_917_out;
            end
        end
        
        assign out_data[917] = lut_917_ff;
    end
    else begin : no_ff_917
        assign out_data[917] = lut_917_out;
    end
    endgenerate
    
    
    
    // LUT : 918
    wire [15:0] lut_918_table = 16'b1100110011110001;
    wire [3:0] lut_918_select = {
                             in_data[154],
                             in_data[424],
                             in_data[209],
                             in_data[556]};
    
    wire lut_918_out = lut_918_table[lut_918_select];
    
    generate
    if ( USE_REG ) begin : ff_918
        reg   lut_918_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_918_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_918_ff <= lut_918_out;
            end
        end
        
        assign out_data[918] = lut_918_ff;
    end
    else begin : no_ff_918
        assign out_data[918] = lut_918_out;
    end
    endgenerate
    
    
    
    // LUT : 919
    wire [15:0] lut_919_table = 16'b1111000111001100;
    wire [3:0] lut_919_select = {
                             in_data[567],
                             in_data[681],
                             in_data[579],
                             in_data[717]};
    
    wire lut_919_out = lut_919_table[lut_919_select];
    
    generate
    if ( USE_REG ) begin : ff_919
        reg   lut_919_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_919_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_919_ff <= lut_919_out;
            end
        end
        
        assign out_data[919] = lut_919_ff;
    end
    else begin : no_ff_919
        assign out_data[919] = lut_919_out;
    end
    endgenerate
    
    
    
    // LUT : 920
    wire [15:0] lut_920_table = 16'b1110111001110111;
    wire [3:0] lut_920_select = {
                             in_data[237],
                             in_data[669],
                             in_data[541],
                             in_data[432]};
    
    wire lut_920_out = lut_920_table[lut_920_select];
    
    generate
    if ( USE_REG ) begin : ff_920
        reg   lut_920_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_920_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_920_ff <= lut_920_out;
            end
        end
        
        assign out_data[920] = lut_920_ff;
    end
    else begin : no_ff_920
        assign out_data[920] = lut_920_out;
    end
    endgenerate
    
    
    
    // LUT : 921
    wire [15:0] lut_921_table = 16'b0001000100010001;
    wire [3:0] lut_921_select = {
                             in_data[645],
                             in_data[23],
                             in_data[479],
                             in_data[245]};
    
    wire lut_921_out = lut_921_table[lut_921_select];
    
    generate
    if ( USE_REG ) begin : ff_921
        reg   lut_921_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_921_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_921_ff <= lut_921_out;
            end
        end
        
        assign out_data[921] = lut_921_ff;
    end
    else begin : no_ff_921
        assign out_data[921] = lut_921_out;
    end
    endgenerate
    
    
    
    // LUT : 922
    wire [15:0] lut_922_table = 16'b1111111110101010;
    wire [3:0] lut_922_select = {
                             in_data[769],
                             in_data[25],
                             in_data[757],
                             in_data[778]};
    
    wire lut_922_out = lut_922_table[lut_922_select];
    
    generate
    if ( USE_REG ) begin : ff_922
        reg   lut_922_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_922_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_922_ff <= lut_922_out;
            end
        end
        
        assign out_data[922] = lut_922_ff;
    end
    else begin : no_ff_922
        assign out_data[922] = lut_922_out;
    end
    endgenerate
    
    
    
    // LUT : 923
    wire [15:0] lut_923_table = 16'b1111111111101110;
    wire [3:0] lut_923_select = {
                             in_data[553],
                             in_data[646],
                             in_data[654],
                             in_data[118]};
    
    wire lut_923_out = lut_923_table[lut_923_select];
    
    generate
    if ( USE_REG ) begin : ff_923
        reg   lut_923_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_923_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_923_ff <= lut_923_out;
            end
        end
        
        assign out_data[923] = lut_923_ff;
    end
    else begin : no_ff_923
        assign out_data[923] = lut_923_out;
    end
    endgenerate
    
    
    
    // LUT : 924
    wire [15:0] lut_924_table = 16'b0000000100000001;
    wire [3:0] lut_924_select = {
                             in_data[5],
                             in_data[201],
                             in_data[98],
                             in_data[147]};
    
    wire lut_924_out = lut_924_table[lut_924_select];
    
    generate
    if ( USE_REG ) begin : ff_924
        reg   lut_924_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_924_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_924_ff <= lut_924_out;
            end
        end
        
        assign out_data[924] = lut_924_ff;
    end
    else begin : no_ff_924
        assign out_data[924] = lut_924_out;
    end
    endgenerate
    
    
    
    // LUT : 925
    wire [15:0] lut_925_table = 16'b1000100011011101;
    wire [3:0] lut_925_select = {
                             in_data[667],
                             in_data[760],
                             in_data[773],
                             in_data[380]};
    
    wire lut_925_out = lut_925_table[lut_925_select];
    
    generate
    if ( USE_REG ) begin : ff_925
        reg   lut_925_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_925_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_925_ff <= lut_925_out;
            end
        end
        
        assign out_data[925] = lut_925_ff;
    end
    else begin : no_ff_925
        assign out_data[925] = lut_925_out;
    end
    endgenerate
    
    
    
    // LUT : 926
    wire [15:0] lut_926_table = 16'b0000001100000011;
    wire [3:0] lut_926_select = {
                             in_data[762],
                             in_data[124],
                             in_data[101],
                             in_data[189]};
    
    wire lut_926_out = lut_926_table[lut_926_select];
    
    generate
    if ( USE_REG ) begin : ff_926
        reg   lut_926_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_926_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_926_ff <= lut_926_out;
            end
        end
        
        assign out_data[926] = lut_926_ff;
    end
    else begin : no_ff_926
        assign out_data[926] = lut_926_out;
    end
    endgenerate
    
    
    
    // LUT : 927
    wire [15:0] lut_927_table = 16'b1111111111110011;
    wire [3:0] lut_927_select = {
                             in_data[355],
                             in_data[302],
                             in_data[519],
                             in_data[722]};
    
    wire lut_927_out = lut_927_table[lut_927_select];
    
    generate
    if ( USE_REG ) begin : ff_927
        reg   lut_927_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_927_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_927_ff <= lut_927_out;
            end
        end
        
        assign out_data[927] = lut_927_ff;
    end
    else begin : no_ff_927
        assign out_data[927] = lut_927_out;
    end
    endgenerate
    
    
    
    // LUT : 928
    wire [15:0] lut_928_table = 16'b0011000011111101;
    wire [3:0] lut_928_select = {
                             in_data[323],
                             in_data[608],
                             in_data[410],
                             in_data[280]};
    
    wire lut_928_out = lut_928_table[lut_928_select];
    
    generate
    if ( USE_REG ) begin : ff_928
        reg   lut_928_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_928_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_928_ff <= lut_928_out;
            end
        end
        
        assign out_data[928] = lut_928_ff;
    end
    else begin : no_ff_928
        assign out_data[928] = lut_928_out;
    end
    endgenerate
    
    
    
    // LUT : 929
    wire [15:0] lut_929_table = 16'b0011111100001001;
    wire [3:0] lut_929_select = {
                             in_data[435],
                             in_data[211],
                             in_data[262],
                             in_data[115]};
    
    wire lut_929_out = lut_929_table[lut_929_select];
    
    generate
    if ( USE_REG ) begin : ff_929
        reg   lut_929_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_929_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_929_ff <= lut_929_out;
            end
        end
        
        assign out_data[929] = lut_929_ff;
    end
    else begin : no_ff_929
        assign out_data[929] = lut_929_out;
    end
    endgenerate
    
    
    
    // LUT : 930
    wire [15:0] lut_930_table = 16'b1000111100001010;
    wire [3:0] lut_930_select = {
                             in_data[507],
                             in_data[482],
                             in_data[412],
                             in_data[293]};
    
    wire lut_930_out = lut_930_table[lut_930_select];
    
    generate
    if ( USE_REG ) begin : ff_930
        reg   lut_930_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_930_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_930_ff <= lut_930_out;
            end
        end
        
        assign out_data[930] = lut_930_ff;
    end
    else begin : no_ff_930
        assign out_data[930] = lut_930_out;
    end
    endgenerate
    
    
    
    // LUT : 931
    wire [15:0] lut_931_table = 16'b0000001000000101;
    wire [3:0] lut_931_select = {
                             in_data[495],
                             in_data[637],
                             in_data[58],
                             in_data[71]};
    
    wire lut_931_out = lut_931_table[lut_931_select];
    
    generate
    if ( USE_REG ) begin : ff_931
        reg   lut_931_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_931_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_931_ff <= lut_931_out;
            end
        end
        
        assign out_data[931] = lut_931_ff;
    end
    else begin : no_ff_931
        assign out_data[931] = lut_931_out;
    end
    endgenerate
    
    
    
    // LUT : 932
    wire [15:0] lut_932_table = 16'b0010001000110011;
    wire [3:0] lut_932_select = {
                             in_data[527],
                             in_data[703],
                             in_data[184],
                             in_data[547]};
    
    wire lut_932_out = lut_932_table[lut_932_select];
    
    generate
    if ( USE_REG ) begin : ff_932
        reg   lut_932_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_932_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_932_ff <= lut_932_out;
            end
        end
        
        assign out_data[932] = lut_932_ff;
    end
    else begin : no_ff_932
        assign out_data[932] = lut_932_out;
    end
    endgenerate
    
    
    
    // LUT : 933
    wire [15:0] lut_933_table = 16'b0101010011110111;
    wire [3:0] lut_933_select = {
                             in_data[238],
                             in_data[441],
                             in_data[515],
                             in_data[712]};
    
    wire lut_933_out = lut_933_table[lut_933_select];
    
    generate
    if ( USE_REG ) begin : ff_933
        reg   lut_933_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_933_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_933_ff <= lut_933_out;
            end
        end
        
        assign out_data[933] = lut_933_ff;
    end
    else begin : no_ff_933
        assign out_data[933] = lut_933_out;
    end
    endgenerate
    
    
    
    // LUT : 934
    wire [15:0] lut_934_table = 16'b0101000011111111;
    wire [3:0] lut_934_select = {
                             in_data[292],
                             in_data[362],
                             in_data[223],
                             in_data[174]};
    
    wire lut_934_out = lut_934_table[lut_934_select];
    
    generate
    if ( USE_REG ) begin : ff_934
        reg   lut_934_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_934_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_934_ff <= lut_934_out;
            end
        end
        
        assign out_data[934] = lut_934_ff;
    end
    else begin : no_ff_934
        assign out_data[934] = lut_934_out;
    end
    endgenerate
    
    
    
    // LUT : 935
    wire [15:0] lut_935_table = 16'b1111111111110000;
    wire [3:0] lut_935_select = {
                             in_data[684],
                             in_data[675],
                             in_data[725],
                             in_data[20]};
    
    wire lut_935_out = lut_935_table[lut_935_select];
    
    generate
    if ( USE_REG ) begin : ff_935
        reg   lut_935_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_935_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_935_ff <= lut_935_out;
            end
        end
        
        assign out_data[935] = lut_935_ff;
    end
    else begin : no_ff_935
        assign out_data[935] = lut_935_out;
    end
    endgenerate
    
    
    
    // LUT : 936
    wire [15:0] lut_936_table = 16'b1111110111111101;
    wire [3:0] lut_936_select = {
                             in_data[140],
                             in_data[445],
                             in_data[46],
                             in_data[753]};
    
    wire lut_936_out = lut_936_table[lut_936_select];
    
    generate
    if ( USE_REG ) begin : ff_936
        reg   lut_936_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_936_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_936_ff <= lut_936_out;
            end
        end
        
        assign out_data[936] = lut_936_ff;
    end
    else begin : no_ff_936
        assign out_data[936] = lut_936_out;
    end
    endgenerate
    
    
    
    // LUT : 937
    wire [15:0] lut_937_table = 16'b1011101110111011;
    wire [3:0] lut_937_select = {
                             in_data[8],
                             in_data[531],
                             in_data[351],
                             in_data[260]};
    
    wire lut_937_out = lut_937_table[lut_937_select];
    
    generate
    if ( USE_REG ) begin : ff_937
        reg   lut_937_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_937_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_937_ff <= lut_937_out;
            end
        end
        
        assign out_data[937] = lut_937_ff;
    end
    else begin : no_ff_937
        assign out_data[937] = lut_937_out;
    end
    endgenerate
    
    
    
    // LUT : 938
    wire [15:0] lut_938_table = 16'b0000001000100011;
    wire [3:0] lut_938_select = {
                             in_data[340],
                             in_data[236],
                             in_data[770],
                             in_data[430]};
    
    wire lut_938_out = lut_938_table[lut_938_select];
    
    generate
    if ( USE_REG ) begin : ff_938
        reg   lut_938_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_938_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_938_ff <= lut_938_out;
            end
        end
        
        assign out_data[938] = lut_938_ff;
    end
    else begin : no_ff_938
        assign out_data[938] = lut_938_out;
    end
    endgenerate
    
    
    
    // LUT : 939
    wire [15:0] lut_939_table = 16'b1111111011111010;
    wire [3:0] lut_939_select = {
                             in_data[192],
                             in_data[374],
                             in_data[549],
                             in_data[613]};
    
    wire lut_939_out = lut_939_table[lut_939_select];
    
    generate
    if ( USE_REG ) begin : ff_939
        reg   lut_939_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_939_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_939_ff <= lut_939_out;
            end
        end
        
        assign out_data[939] = lut_939_ff;
    end
    else begin : no_ff_939
        assign out_data[939] = lut_939_out;
    end
    endgenerate
    
    
    
    // LUT : 940
    wire [15:0] lut_940_table = 16'b1111111111111101;
    wire [3:0] lut_940_select = {
                             in_data[171],
                             in_data[77],
                             in_data[529],
                             in_data[31]};
    
    wire lut_940_out = lut_940_table[lut_940_select];
    
    generate
    if ( USE_REG ) begin : ff_940
        reg   lut_940_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_940_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_940_ff <= lut_940_out;
            end
        end
        
        assign out_data[940] = lut_940_ff;
    end
    else begin : no_ff_940
        assign out_data[940] = lut_940_out;
    end
    endgenerate
    
    
    
    // LUT : 941
    wire [15:0] lut_941_table = 16'b0000000011111111;
    wire [3:0] lut_941_select = {
                             in_data[409],
                             in_data[642],
                             in_data[213],
                             in_data[369]};
    
    wire lut_941_out = lut_941_table[lut_941_select];
    
    generate
    if ( USE_REG ) begin : ff_941
        reg   lut_941_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_941_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_941_ff <= lut_941_out;
            end
        end
        
        assign out_data[941] = lut_941_ff;
    end
    else begin : no_ff_941
        assign out_data[941] = lut_941_out;
    end
    endgenerate
    
    
    
    // LUT : 942
    wire [15:0] lut_942_table = 16'b0000000000000011;
    wire [3:0] lut_942_select = {
                             in_data[386],
                             in_data[464],
                             in_data[457],
                             in_data[700]};
    
    wire lut_942_out = lut_942_table[lut_942_select];
    
    generate
    if ( USE_REG ) begin : ff_942
        reg   lut_942_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_942_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_942_ff <= lut_942_out;
            end
        end
        
        assign out_data[942] = lut_942_ff;
    end
    else begin : no_ff_942
        assign out_data[942] = lut_942_out;
    end
    endgenerate
    
    
    
    // LUT : 943
    wire [15:0] lut_943_table = 16'b0000001000000010;
    wire [3:0] lut_943_select = {
                             in_data[782],
                             in_data[277],
                             in_data[250],
                             in_data[520]};
    
    wire lut_943_out = lut_943_table[lut_943_select];
    
    generate
    if ( USE_REG ) begin : ff_943
        reg   lut_943_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_943_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_943_ff <= lut_943_out;
            end
        end
        
        assign out_data[943] = lut_943_ff;
    end
    else begin : no_ff_943
        assign out_data[943] = lut_943_out;
    end
    endgenerate
    
    
    
    // LUT : 944
    wire [15:0] lut_944_table = 16'b0000111000000011;
    wire [3:0] lut_944_select = {
                             in_data[347],
                             in_data[639],
                             in_data[148],
                             in_data[389]};
    
    wire lut_944_out = lut_944_table[lut_944_select];
    
    generate
    if ( USE_REG ) begin : ff_944
        reg   lut_944_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_944_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_944_ff <= lut_944_out;
            end
        end
        
        assign out_data[944] = lut_944_ff;
    end
    else begin : no_ff_944
        assign out_data[944] = lut_944_out;
    end
    endgenerate
    
    
    
    // LUT : 945
    wire [15:0] lut_945_table = 16'b0000000000000101;
    wire [3:0] lut_945_select = {
                             in_data[473],
                             in_data[281],
                             in_data[4],
                             in_data[413]};
    
    wire lut_945_out = lut_945_table[lut_945_select];
    
    generate
    if ( USE_REG ) begin : ff_945
        reg   lut_945_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_945_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_945_ff <= lut_945_out;
            end
        end
        
        assign out_data[945] = lut_945_ff;
    end
    else begin : no_ff_945
        assign out_data[945] = lut_945_out;
    end
    endgenerate
    
    
    
    // LUT : 946
    wire [15:0] lut_946_table = 16'b1111111111001100;
    wire [3:0] lut_946_select = {
                             in_data[568],
                             in_data[224],
                             in_data[650],
                             in_data[755]};
    
    wire lut_946_out = lut_946_table[lut_946_select];
    
    generate
    if ( USE_REG ) begin : ff_946
        reg   lut_946_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_946_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_946_ff <= lut_946_out;
            end
        end
        
        assign out_data[946] = lut_946_ff;
    end
    else begin : no_ff_946
        assign out_data[946] = lut_946_out;
    end
    endgenerate
    
    
    
    // LUT : 947
    wire [15:0] lut_947_table = 16'b1111111111111010;
    wire [3:0] lut_947_select = {
                             in_data[402],
                             in_data[248],
                             in_data[469],
                             in_data[68]};
    
    wire lut_947_out = lut_947_table[lut_947_select];
    
    generate
    if ( USE_REG ) begin : ff_947
        reg   lut_947_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_947_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_947_ff <= lut_947_out;
            end
        end
        
        assign out_data[947] = lut_947_ff;
    end
    else begin : no_ff_947
        assign out_data[947] = lut_947_out;
    end
    endgenerate
    
    
    
    // LUT : 948
    wire [15:0] lut_948_table = 16'b1111111011101110;
    wire [3:0] lut_948_select = {
                             in_data[233],
                             in_data[273],
                             in_data[737],
                             in_data[379]};
    
    wire lut_948_out = lut_948_table[lut_948_select];
    
    generate
    if ( USE_REG ) begin : ff_948
        reg   lut_948_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_948_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_948_ff <= lut_948_out;
            end
        end
        
        assign out_data[948] = lut_948_ff;
    end
    else begin : no_ff_948
        assign out_data[948] = lut_948_out;
    end
    endgenerate
    
    
    
    // LUT : 949
    wire [15:0] lut_949_table = 16'b1111101100110010;
    wire [3:0] lut_949_select = {
                             in_data[221],
                             in_data[396],
                             in_data[648],
                             in_data[750]};
    
    wire lut_949_out = lut_949_table[lut_949_select];
    
    generate
    if ( USE_REG ) begin : ff_949
        reg   lut_949_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_949_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_949_ff <= lut_949_out;
            end
        end
        
        assign out_data[949] = lut_949_ff;
    end
    else begin : no_ff_949
        assign out_data[949] = lut_949_out;
    end
    endgenerate
    
    
    
    // LUT : 950
    wire [15:0] lut_950_table = 16'b0000110101001101;
    wire [3:0] lut_950_select = {
                             in_data[443],
                             in_data[427],
                             in_data[744],
                             in_data[160]};
    
    wire lut_950_out = lut_950_table[lut_950_select];
    
    generate
    if ( USE_REG ) begin : ff_950
        reg   lut_950_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_950_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_950_ff <= lut_950_out;
            end
        end
        
        assign out_data[950] = lut_950_ff;
    end
    else begin : no_ff_950
        assign out_data[950] = lut_950_out;
    end
    endgenerate
    
    
    
    // LUT : 951
    wire [15:0] lut_951_table = 16'b1111111111111110;
    wire [3:0] lut_951_select = {
                             in_data[228],
                             in_data[338],
                             in_data[332],
                             in_data[377]};
    
    wire lut_951_out = lut_951_table[lut_951_select];
    
    generate
    if ( USE_REG ) begin : ff_951
        reg   lut_951_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_951_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_951_ff <= lut_951_out;
            end
        end
        
        assign out_data[951] = lut_951_ff;
    end
    else begin : no_ff_951
        assign out_data[951] = lut_951_out;
    end
    endgenerate
    
    
    
    // LUT : 952
    wire [15:0] lut_952_table = 16'b1000000000100010;
    wire [3:0] lut_952_select = {
                             in_data[584],
                             in_data[127],
                             in_data[581],
                             in_data[300]};
    
    wire lut_952_out = lut_952_table[lut_952_select];
    
    generate
    if ( USE_REG ) begin : ff_952
        reg   lut_952_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_952_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_952_ff <= lut_952_out;
            end
        end
        
        assign out_data[952] = lut_952_ff;
    end
    else begin : no_ff_952
        assign out_data[952] = lut_952_out;
    end
    endgenerate
    
    
    
    // LUT : 953
    wire [15:0] lut_953_table = 16'b1111111100000000;
    wire [3:0] lut_953_select = {
                             in_data[301],
                             in_data[638],
                             in_data[196],
                             in_data[510]};
    
    wire lut_953_out = lut_953_table[lut_953_select];
    
    generate
    if ( USE_REG ) begin : ff_953
        reg   lut_953_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_953_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_953_ff <= lut_953_out;
            end
        end
        
        assign out_data[953] = lut_953_ff;
    end
    else begin : no_ff_953
        assign out_data[953] = lut_953_out;
    end
    endgenerate
    
    
    
    // LUT : 954
    wire [15:0] lut_954_table = 16'b0100010100000101;
    wire [3:0] lut_954_select = {
                             in_data[502],
                             in_data[134],
                             in_data[282],
                             in_data[247]};
    
    wire lut_954_out = lut_954_table[lut_954_select];
    
    generate
    if ( USE_REG ) begin : ff_954
        reg   lut_954_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_954_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_954_ff <= lut_954_out;
            end
        end
        
        assign out_data[954] = lut_954_ff;
    end
    else begin : no_ff_954
        assign out_data[954] = lut_954_out;
    end
    endgenerate
    
    
    
    // LUT : 955
    wire [15:0] lut_955_table = 16'b1111111111111010;
    wire [3:0] lut_955_select = {
                             in_data[752],
                             in_data[60],
                             in_data[56],
                             in_data[202]};
    
    wire lut_955_out = lut_955_table[lut_955_select];
    
    generate
    if ( USE_REG ) begin : ff_955
        reg   lut_955_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_955_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_955_ff <= lut_955_out;
            end
        end
        
        assign out_data[955] = lut_955_ff;
    end
    else begin : no_ff_955
        assign out_data[955] = lut_955_out;
    end
    endgenerate
    
    
    
    // LUT : 956
    wire [15:0] lut_956_table = 16'b1111111111001100;
    wire [3:0] lut_956_select = {
                             in_data[632],
                             in_data[286],
                             in_data[107],
                             in_data[3]};
    
    wire lut_956_out = lut_956_table[lut_956_select];
    
    generate
    if ( USE_REG ) begin : ff_956
        reg   lut_956_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_956_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_956_ff <= lut_956_out;
            end
        end
        
        assign out_data[956] = lut_956_ff;
    end
    else begin : no_ff_956
        assign out_data[956] = lut_956_out;
    end
    endgenerate
    
    
    
    // LUT : 957
    wire [15:0] lut_957_table = 16'b1111111111011101;
    wire [3:0] lut_957_select = {
                             in_data[511],
                             in_data[320],
                             in_data[246],
                             in_data[182]};
    
    wire lut_957_out = lut_957_table[lut_957_select];
    
    generate
    if ( USE_REG ) begin : ff_957
        reg   lut_957_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_957_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_957_ff <= lut_957_out;
            end
        end
        
        assign out_data[957] = lut_957_ff;
    end
    else begin : no_ff_957
        assign out_data[957] = lut_957_out;
    end
    endgenerate
    
    
    
    // LUT : 958
    wire [15:0] lut_958_table = 16'b1010101011111010;
    wire [3:0] lut_958_select = {
                             in_data[429],
                             in_data[434],
                             in_data[49],
                             in_data[311]};
    
    wire lut_958_out = lut_958_table[lut_958_select];
    
    generate
    if ( USE_REG ) begin : ff_958
        reg   lut_958_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_958_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_958_ff <= lut_958_out;
            end
        end
        
        assign out_data[958] = lut_958_ff;
    end
    else begin : no_ff_958
        assign out_data[958] = lut_958_out;
    end
    endgenerate
    
    
    
    // LUT : 959
    wire [15:0] lut_959_table = 16'b1000100010001100;
    wire [3:0] lut_959_select = {
                             in_data[401],
                             in_data[569],
                             in_data[269],
                             in_data[378]};
    
    wire lut_959_out = lut_959_table[lut_959_select];
    
    generate
    if ( USE_REG ) begin : ff_959
        reg   lut_959_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_959_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_959_ff <= lut_959_out;
            end
        end
        
        assign out_data[959] = lut_959_ff;
    end
    else begin : no_ff_959
        assign out_data[959] = lut_959_out;
    end
    endgenerate
    
    
    
    // LUT : 960
    wire [15:0] lut_960_table = 16'b1111001111110000;
    wire [3:0] lut_960_select = {
                             in_data[244],
                             in_data[229],
                             in_data[249],
                             in_data[698]};
    
    wire lut_960_out = lut_960_table[lut_960_select];
    
    generate
    if ( USE_REG ) begin : ff_960
        reg   lut_960_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_960_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_960_ff <= lut_960_out;
            end
        end
        
        assign out_data[960] = lut_960_ff;
    end
    else begin : no_ff_960
        assign out_data[960] = lut_960_out;
    end
    endgenerate
    
    
    
    // LUT : 961
    wire [15:0] lut_961_table = 16'b0000000001111100;
    wire [3:0] lut_961_select = {
                             in_data[562],
                             in_data[664],
                             in_data[318],
                             in_data[641]};
    
    wire lut_961_out = lut_961_table[lut_961_select];
    
    generate
    if ( USE_REG ) begin : ff_961
        reg   lut_961_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_961_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_961_ff <= lut_961_out;
            end
        end
        
        assign out_data[961] = lut_961_ff;
    end
    else begin : no_ff_961
        assign out_data[961] = lut_961_out;
    end
    endgenerate
    
    
    
    // LUT : 962
    wire [15:0] lut_962_table = 16'b0010001011111111;
    wire [3:0] lut_962_select = {
                             in_data[517],
                             in_data[16],
                             in_data[509],
                             in_data[305]};
    
    wire lut_962_out = lut_962_table[lut_962_select];
    
    generate
    if ( USE_REG ) begin : ff_962
        reg   lut_962_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_962_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_962_ff <= lut_962_out;
            end
        end
        
        assign out_data[962] = lut_962_ff;
    end
    else begin : no_ff_962
        assign out_data[962] = lut_962_out;
    end
    endgenerate
    
    
    
    // LUT : 963
    wire [15:0] lut_963_table = 16'b1111111111111110;
    wire [3:0] lut_963_select = {
                             in_data[131],
                             in_data[720],
                             in_data[162],
                             in_data[694]};
    
    wire lut_963_out = lut_963_table[lut_963_select];
    
    generate
    if ( USE_REG ) begin : ff_963
        reg   lut_963_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_963_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_963_ff <= lut_963_out;
            end
        end
        
        assign out_data[963] = lut_963_ff;
    end
    else begin : no_ff_963
        assign out_data[963] = lut_963_out;
    end
    endgenerate
    
    
    
    // LUT : 964
    wire [15:0] lut_964_table = 16'b1101111100000000;
    wire [3:0] lut_964_select = {
                             in_data[316],
                             in_data[595],
                             in_data[258],
                             in_data[601]};
    
    wire lut_964_out = lut_964_table[lut_964_select];
    
    generate
    if ( USE_REG ) begin : ff_964
        reg   lut_964_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_964_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_964_ff <= lut_964_out;
            end
        end
        
        assign out_data[964] = lut_964_ff;
    end
    else begin : no_ff_964
        assign out_data[964] = lut_964_out;
    end
    endgenerate
    
    
    
    // LUT : 965
    wire [15:0] lut_965_table = 16'b0000000100000001;
    wire [3:0] lut_965_select = {
                             in_data[578],
                             in_data[506],
                             in_data[296],
                             in_data[706]};
    
    wire lut_965_out = lut_965_table[lut_965_select];
    
    generate
    if ( USE_REG ) begin : ff_965
        reg   lut_965_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_965_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_965_ff <= lut_965_out;
            end
        end
        
        assign out_data[965] = lut_965_ff;
    end
    else begin : no_ff_965
        assign out_data[965] = lut_965_out;
    end
    endgenerate
    
    
    
    // LUT : 966
    wire [15:0] lut_966_table = 16'b1111111011001100;
    wire [3:0] lut_966_select = {
                             in_data[69],
                             in_data[551],
                             in_data[235],
                             in_data[746]};
    
    wire lut_966_out = lut_966_table[lut_966_select];
    
    generate
    if ( USE_REG ) begin : ff_966
        reg   lut_966_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_966_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_966_ff <= lut_966_out;
            end
        end
        
        assign out_data[966] = lut_966_ff;
    end
    else begin : no_ff_966
        assign out_data[966] = lut_966_out;
    end
    endgenerate
    
    
    
    // LUT : 967
    wire [15:0] lut_967_table = 16'b1111000011110000;
    wire [3:0] lut_967_select = {
                             in_data[392],
                             in_data[518],
                             in_data[423],
                             in_data[38]};
    
    wire lut_967_out = lut_967_table[lut_967_select];
    
    generate
    if ( USE_REG ) begin : ff_967
        reg   lut_967_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_967_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_967_ff <= lut_967_out;
            end
        end
        
        assign out_data[967] = lut_967_ff;
    end
    else begin : no_ff_967
        assign out_data[967] = lut_967_out;
    end
    endgenerate
    
    
    
    // LUT : 968
    wire [15:0] lut_968_table = 16'b1111111111101110;
    wire [3:0] lut_968_select = {
                             in_data[481],
                             in_data[604],
                             in_data[439],
                             in_data[400]};
    
    wire lut_968_out = lut_968_table[lut_968_select];
    
    generate
    if ( USE_REG ) begin : ff_968
        reg   lut_968_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_968_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_968_ff <= lut_968_out;
            end
        end
        
        assign out_data[968] = lut_968_ff;
    end
    else begin : no_ff_968
        assign out_data[968] = lut_968_out;
    end
    endgenerate
    
    
    
    // LUT : 969
    wire [15:0] lut_969_table = 16'b0000000000001110;
    wire [3:0] lut_969_select = {
                             in_data[255],
                             in_data[539],
                             in_data[468],
                             in_data[612]};
    
    wire lut_969_out = lut_969_table[lut_969_select];
    
    generate
    if ( USE_REG ) begin : ff_969
        reg   lut_969_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_969_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_969_ff <= lut_969_out;
            end
        end
        
        assign out_data[969] = lut_969_ff;
    end
    else begin : no_ff_969
        assign out_data[969] = lut_969_out;
    end
    endgenerate
    
    
    
    // LUT : 970
    wire [15:0] lut_970_table = 16'b0101010100010001;
    wire [3:0] lut_970_select = {
                             in_data[366],
                             in_data[2],
                             in_data[90],
                             in_data[122]};
    
    wire lut_970_out = lut_970_table[lut_970_select];
    
    generate
    if ( USE_REG ) begin : ff_970
        reg   lut_970_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_970_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_970_ff <= lut_970_out;
            end
        end
        
        assign out_data[970] = lut_970_ff;
    end
    else begin : no_ff_970
        assign out_data[970] = lut_970_out;
    end
    endgenerate
    
    
    
    // LUT : 971
    wire [15:0] lut_971_table = 16'b0011001100010000;
    wire [3:0] lut_971_select = {
                             in_data[690],
                             in_data[34],
                             in_data[120],
                             in_data[226]};
    
    wire lut_971_out = lut_971_table[lut_971_select];
    
    generate
    if ( USE_REG ) begin : ff_971
        reg   lut_971_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_971_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_971_ff <= lut_971_out;
            end
        end
        
        assign out_data[971] = lut_971_ff;
    end
    else begin : no_ff_971
        assign out_data[971] = lut_971_out;
    end
    endgenerate
    
    
    
    // LUT : 972
    wire [15:0] lut_972_table = 16'b1010111100001111;
    wire [3:0] lut_972_select = {
                             in_data[484],
                             in_data[267],
                             in_data[337],
                             in_data[723]};
    
    wire lut_972_out = lut_972_table[lut_972_select];
    
    generate
    if ( USE_REG ) begin : ff_972
        reg   lut_972_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_972_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_972_ff <= lut_972_out;
            end
        end
        
        assign out_data[972] = lut_972_ff;
    end
    else begin : no_ff_972
        assign out_data[972] = lut_972_out;
    end
    endgenerate
    
    
    
    // LUT : 973
    wire [15:0] lut_973_table = 16'b0000000000000011;
    wire [3:0] lut_973_select = {
                             in_data[283],
                             in_data[425],
                             in_data[523],
                             in_data[749]};
    
    wire lut_973_out = lut_973_table[lut_973_select];
    
    generate
    if ( USE_REG ) begin : ff_973
        reg   lut_973_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_973_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_973_ff <= lut_973_out;
            end
        end
        
        assign out_data[973] = lut_973_ff;
    end
    else begin : no_ff_973
        assign out_data[973] = lut_973_out;
    end
    endgenerate
    
    
    
    // LUT : 974
    wire [15:0] lut_974_table = 16'b1011001010100011;
    wire [3:0] lut_974_select = {
                             in_data[290],
                             in_data[415],
                             in_data[289],
                             in_data[704]};
    
    wire lut_974_out = lut_974_table[lut_974_select];
    
    generate
    if ( USE_REG ) begin : ff_974
        reg   lut_974_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_974_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_974_ff <= lut_974_out;
            end
        end
        
        assign out_data[974] = lut_974_ff;
    end
    else begin : no_ff_974
        assign out_data[974] = lut_974_out;
    end
    endgenerate
    
    
    
    // LUT : 975
    wire [15:0] lut_975_table = 16'b0000000000001111;
    wire [3:0] lut_975_select = {
                             in_data[136],
                             in_data[313],
                             in_data[751],
                             in_data[117]};
    
    wire lut_975_out = lut_975_table[lut_975_select];
    
    generate
    if ( USE_REG ) begin : ff_975
        reg   lut_975_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_975_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_975_ff <= lut_975_out;
            end
        end
        
        assign out_data[975] = lut_975_ff;
    end
    else begin : no_ff_975
        assign out_data[975] = lut_975_out;
    end
    endgenerate
    
    
    
    // LUT : 976
    wire [15:0] lut_976_table = 16'b1111111111111110;
    wire [3:0] lut_976_select = {
                             in_data[252],
                             in_data[55],
                             in_data[50],
                             in_data[677]};
    
    wire lut_976_out = lut_976_table[lut_976_select];
    
    generate
    if ( USE_REG ) begin : ff_976
        reg   lut_976_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_976_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_976_ff <= lut_976_out;
            end
        end
        
        assign out_data[976] = lut_976_ff;
    end
    else begin : no_ff_976
        assign out_data[976] = lut_976_out;
    end
    endgenerate
    
    
    
    // LUT : 977
    wire [15:0] lut_977_table = 16'b1011101010111110;
    wire [3:0] lut_977_select = {
                             in_data[580],
                             in_data[453],
                             in_data[385],
                             in_data[598]};
    
    wire lut_977_out = lut_977_table[lut_977_select];
    
    generate
    if ( USE_REG ) begin : ff_977
        reg   lut_977_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_977_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_977_ff <= lut_977_out;
            end
        end
        
        assign out_data[977] = lut_977_ff;
    end
    else begin : no_ff_977
        assign out_data[977] = lut_977_out;
    end
    endgenerate
    
    
    
    // LUT : 978
    wire [15:0] lut_978_table = 16'b1111101111010011;
    wire [3:0] lut_978_select = {
                             in_data[411],
                             in_data[653],
                             in_data[266],
                             in_data[241]};
    
    wire lut_978_out = lut_978_table[lut_978_select];
    
    generate
    if ( USE_REG ) begin : ff_978
        reg   lut_978_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_978_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_978_ff <= lut_978_out;
            end
        end
        
        assign out_data[978] = lut_978_ff;
    end
    else begin : no_ff_978
        assign out_data[978] = lut_978_out;
    end
    endgenerate
    
    
    
    // LUT : 979
    wire [15:0] lut_979_table = 16'b0010101010101011;
    wire [3:0] lut_979_select = {
                             in_data[76],
                             in_data[573],
                             in_data[130],
                             in_data[661]};
    
    wire lut_979_out = lut_979_table[lut_979_select];
    
    generate
    if ( USE_REG ) begin : ff_979
        reg   lut_979_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_979_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_979_ff <= lut_979_out;
            end
        end
        
        assign out_data[979] = lut_979_ff;
    end
    else begin : no_ff_979
        assign out_data[979] = lut_979_out;
    end
    endgenerate
    
    
    
    // LUT : 980
    wire [15:0] lut_980_table = 16'b1111000011111110;
    wire [3:0] lut_980_select = {
                             in_data[258],
                             in_data[548],
                             in_data[618],
                             in_data[441]};
    
    wire lut_980_out = lut_980_table[lut_980_select];
    
    generate
    if ( USE_REG ) begin : ff_980
        reg   lut_980_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_980_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_980_ff <= lut_980_out;
            end
        end
        
        assign out_data[980] = lut_980_ff;
    end
    else begin : no_ff_980
        assign out_data[980] = lut_980_out;
    end
    endgenerate
    
    
    
    // LUT : 981
    wire [15:0] lut_981_table = 16'b0111000101110001;
    wire [3:0] lut_981_select = {
                             in_data[752],
                             in_data[499],
                             in_data[187],
                             in_data[437]};
    
    wire lut_981_out = lut_981_table[lut_981_select];
    
    generate
    if ( USE_REG ) begin : ff_981
        reg   lut_981_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_981_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_981_ff <= lut_981_out;
            end
        end
        
        assign out_data[981] = lut_981_ff;
    end
    else begin : no_ff_981
        assign out_data[981] = lut_981_out;
    end
    endgenerate
    
    
    
    // LUT : 982
    wire [15:0] lut_982_table = 16'b1111101011111111;
    wire [3:0] lut_982_select = {
                             in_data[463],
                             in_data[277],
                             in_data[617],
                             in_data[412]};
    
    wire lut_982_out = lut_982_table[lut_982_select];
    
    generate
    if ( USE_REG ) begin : ff_982
        reg   lut_982_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_982_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_982_ff <= lut_982_out;
            end
        end
        
        assign out_data[982] = lut_982_ff;
    end
    else begin : no_ff_982
        assign out_data[982] = lut_982_out;
    end
    endgenerate
    
    
    
    // LUT : 983
    wire [15:0] lut_983_table = 16'b0000000000000101;
    wire [3:0] lut_983_select = {
                             in_data[174],
                             in_data[294],
                             in_data[421],
                             in_data[541]};
    
    wire lut_983_out = lut_983_table[lut_983_select];
    
    generate
    if ( USE_REG ) begin : ff_983
        reg   lut_983_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_983_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_983_ff <= lut_983_out;
            end
        end
        
        assign out_data[983] = lut_983_ff;
    end
    else begin : no_ff_983
        assign out_data[983] = lut_983_out;
    end
    endgenerate
    
    
    
    // LUT : 984
    wire [15:0] lut_984_table = 16'b1111110011111100;
    wire [3:0] lut_984_select = {
                             in_data[338],
                             in_data[605],
                             in_data[557],
                             in_data[59]};
    
    wire lut_984_out = lut_984_table[lut_984_select];
    
    generate
    if ( USE_REG ) begin : ff_984
        reg   lut_984_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_984_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_984_ff <= lut_984_out;
            end
        end
        
        assign out_data[984] = lut_984_ff;
    end
    else begin : no_ff_984
        assign out_data[984] = lut_984_out;
    end
    endgenerate
    
    
    
    // LUT : 985
    wire [15:0] lut_985_table = 16'b0101010101010101;
    wire [3:0] lut_985_select = {
                             in_data[7],
                             in_data[139],
                             in_data[454],
                             in_data[320]};
    
    wire lut_985_out = lut_985_table[lut_985_select];
    
    generate
    if ( USE_REG ) begin : ff_985
        reg   lut_985_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_985_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_985_ff <= lut_985_out;
            end
        end
        
        assign out_data[985] = lut_985_ff;
    end
    else begin : no_ff_985
        assign out_data[985] = lut_985_out;
    end
    endgenerate
    
    
    
    // LUT : 986
    wire [15:0] lut_986_table = 16'b0000000000000001;
    wire [3:0] lut_986_select = {
                             in_data[95],
                             in_data[616],
                             in_data[614],
                             in_data[44]};
    
    wire lut_986_out = lut_986_table[lut_986_select];
    
    generate
    if ( USE_REG ) begin : ff_986
        reg   lut_986_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_986_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_986_ff <= lut_986_out;
            end
        end
        
        assign out_data[986] = lut_986_ff;
    end
    else begin : no_ff_986
        assign out_data[986] = lut_986_out;
    end
    endgenerate
    
    
    
    // LUT : 987
    wire [15:0] lut_987_table = 16'b0000001100000011;
    wire [3:0] lut_987_select = {
                             in_data[698],
                             in_data[691],
                             in_data[265],
                             in_data[264]};
    
    wire lut_987_out = lut_987_table[lut_987_select];
    
    generate
    if ( USE_REG ) begin : ff_987
        reg   lut_987_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_987_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_987_ff <= lut_987_out;
            end
        end
        
        assign out_data[987] = lut_987_ff;
    end
    else begin : no_ff_987
        assign out_data[987] = lut_987_out;
    end
    endgenerate
    
    
    
    // LUT : 988
    wire [15:0] lut_988_table = 16'b0000001100000001;
    wire [3:0] lut_988_select = {
                             in_data[183],
                             in_data[578],
                             in_data[494],
                             in_data[83]};
    
    wire lut_988_out = lut_988_table[lut_988_select];
    
    generate
    if ( USE_REG ) begin : ff_988
        reg   lut_988_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_988_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_988_ff <= lut_988_out;
            end
        end
        
        assign out_data[988] = lut_988_ff;
    end
    else begin : no_ff_988
        assign out_data[988] = lut_988_out;
    end
    endgenerate
    
    
    
    // LUT : 989
    wire [15:0] lut_989_table = 16'b0000000000010001;
    wire [3:0] lut_989_select = {
                             in_data[339],
                             in_data[471],
                             in_data[510],
                             in_data[547]};
    
    wire lut_989_out = lut_989_table[lut_989_select];
    
    generate
    if ( USE_REG ) begin : ff_989
        reg   lut_989_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_989_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_989_ff <= lut_989_out;
            end
        end
        
        assign out_data[989] = lut_989_ff;
    end
    else begin : no_ff_989
        assign out_data[989] = lut_989_out;
    end
    endgenerate
    
    
    
    // LUT : 990
    wire [15:0] lut_990_table = 16'b1111111100000000;
    wire [3:0] lut_990_select = {
                             in_data[376],
                             in_data[117],
                             in_data[28],
                             in_data[478]};
    
    wire lut_990_out = lut_990_table[lut_990_select];
    
    generate
    if ( USE_REG ) begin : ff_990
        reg   lut_990_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_990_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_990_ff <= lut_990_out;
            end
        end
        
        assign out_data[990] = lut_990_ff;
    end
    else begin : no_ff_990
        assign out_data[990] = lut_990_out;
    end
    endgenerate
    
    
    
    // LUT : 991
    wire [15:0] lut_991_table = 16'b0101010100000000;
    wire [3:0] lut_991_select = {
                             in_data[433],
                             in_data[224],
                             in_data[643],
                             in_data[502]};
    
    wire lut_991_out = lut_991_table[lut_991_select];
    
    generate
    if ( USE_REG ) begin : ff_991
        reg   lut_991_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_991_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_991_ff <= lut_991_out;
            end
        end
        
        assign out_data[991] = lut_991_ff;
    end
    else begin : no_ff_991
        assign out_data[991] = lut_991_out;
    end
    endgenerate
    
    
    
    // LUT : 992
    wire [15:0] lut_992_table = 16'b0011001100110011;
    wire [3:0] lut_992_select = {
                             in_data[1],
                             in_data[53],
                             in_data[458],
                             in_data[753]};
    
    wire lut_992_out = lut_992_table[lut_992_select];
    
    generate
    if ( USE_REG ) begin : ff_992
        reg   lut_992_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_992_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_992_ff <= lut_992_out;
            end
        end
        
        assign out_data[992] = lut_992_ff;
    end
    else begin : no_ff_992
        assign out_data[992] = lut_992_out;
    end
    endgenerate
    
    
    
    // LUT : 993
    wire [15:0] lut_993_table = 16'b0100110000001100;
    wire [3:0] lut_993_select = {
                             in_data[130],
                             in_data[746],
                             in_data[426],
                             in_data[118]};
    
    wire lut_993_out = lut_993_table[lut_993_select];
    
    generate
    if ( USE_REG ) begin : ff_993
        reg   lut_993_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_993_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_993_ff <= lut_993_out;
            end
        end
        
        assign out_data[993] = lut_993_ff;
    end
    else begin : no_ff_993
        assign out_data[993] = lut_993_out;
    end
    endgenerate
    
    
    
    // LUT : 994
    wire [15:0] lut_994_table = 16'b0000000011110000;
    wire [3:0] lut_994_select = {
                             in_data[411],
                             in_data[404],
                             in_data[771],
                             in_data[562]};
    
    wire lut_994_out = lut_994_table[lut_994_select];
    
    generate
    if ( USE_REG ) begin : ff_994
        reg   lut_994_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_994_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_994_ff <= lut_994_out;
            end
        end
        
        assign out_data[994] = lut_994_ff;
    end
    else begin : no_ff_994
        assign out_data[994] = lut_994_out;
    end
    endgenerate
    
    
    
    // LUT : 995
    wire [15:0] lut_995_table = 16'b1010111110101010;
    wire [3:0] lut_995_select = {
                             in_data[132],
                             in_data[347],
                             in_data[0],
                             in_data[431]};
    
    wire lut_995_out = lut_995_table[lut_995_select];
    
    generate
    if ( USE_REG ) begin : ff_995
        reg   lut_995_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_995_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_995_ff <= lut_995_out;
            end
        end
        
        assign out_data[995] = lut_995_ff;
    end
    else begin : no_ff_995
        assign out_data[995] = lut_995_out;
    end
    endgenerate
    
    
    
    // LUT : 996
    wire [15:0] lut_996_table = 16'b1111111110101010;
    wire [3:0] lut_996_select = {
                             in_data[739],
                             in_data[631],
                             in_data[507],
                             in_data[343]};
    
    wire lut_996_out = lut_996_table[lut_996_select];
    
    generate
    if ( USE_REG ) begin : ff_996
        reg   lut_996_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_996_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_996_ff <= lut_996_out;
            end
        end
        
        assign out_data[996] = lut_996_ff;
    end
    else begin : no_ff_996
        assign out_data[996] = lut_996_out;
    end
    endgenerate
    
    
    
    // LUT : 997
    wire [15:0] lut_997_table = 16'b1111111111111010;
    wire [3:0] lut_997_select = {
                             in_data[584],
                             in_data[362],
                             in_data[88],
                             in_data[568]};
    
    wire lut_997_out = lut_997_table[lut_997_select];
    
    generate
    if ( USE_REG ) begin : ff_997
        reg   lut_997_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_997_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_997_ff <= lut_997_out;
            end
        end
        
        assign out_data[997] = lut_997_ff;
    end
    else begin : no_ff_997
        assign out_data[997] = lut_997_out;
    end
    endgenerate
    
    
    
    // LUT : 998
    wire [15:0] lut_998_table = 16'b0011111100000011;
    wire [3:0] lut_998_select = {
                             in_data[200],
                             in_data[538],
                             in_data[419],
                             in_data[251]};
    
    wire lut_998_out = lut_998_table[lut_998_select];
    
    generate
    if ( USE_REG ) begin : ff_998
        reg   lut_998_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_998_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_998_ff <= lut_998_out;
            end
        end
        
        assign out_data[998] = lut_998_ff;
    end
    else begin : no_ff_998
        assign out_data[998] = lut_998_out;
    end
    endgenerate
    
    
    
    // LUT : 999
    wire [15:0] lut_999_table = 16'b0000000000000101;
    wire [3:0] lut_999_select = {
                             in_data[255],
                             in_data[274],
                             in_data[18],
                             in_data[748]};
    
    wire lut_999_out = lut_999_table[lut_999_select];
    
    generate
    if ( USE_REG ) begin : ff_999
        reg   lut_999_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_999_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_999_ff <= lut_999_out;
            end
        end
        
        assign out_data[999] = lut_999_ff;
    end
    else begin : no_ff_999
        assign out_data[999] = lut_999_out;
    end
    endgenerate
    
    
    
    // LUT : 1000
    wire [15:0] lut_1000_table = 16'b1111000011111000;
    wire [3:0] lut_1000_select = {
                             in_data[133],
                             in_data[300],
                             in_data[501],
                             in_data[436]};
    
    wire lut_1000_out = lut_1000_table[lut_1000_select];
    
    generate
    if ( USE_REG ) begin : ff_1000
        reg   lut_1000_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1000_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1000_ff <= lut_1000_out;
            end
        end
        
        assign out_data[1000] = lut_1000_ff;
    end
    else begin : no_ff_1000
        assign out_data[1000] = lut_1000_out;
    end
    endgenerate
    
    
    
    // LUT : 1001
    wire [15:0] lut_1001_table = 16'b0000101000001110;
    wire [3:0] lut_1001_select = {
                             in_data[615],
                             in_data[330],
                             in_data[90],
                             in_data[350]};
    
    wire lut_1001_out = lut_1001_table[lut_1001_select];
    
    generate
    if ( USE_REG ) begin : ff_1001
        reg   lut_1001_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1001_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1001_ff <= lut_1001_out;
            end
        end
        
        assign out_data[1001] = lut_1001_ff;
    end
    else begin : no_ff_1001
        assign out_data[1001] = lut_1001_out;
    end
    endgenerate
    
    
    
    // LUT : 1002
    wire [15:0] lut_1002_table = 16'b1111111110110000;
    wire [3:0] lut_1002_select = {
                             in_data[377],
                             in_data[220],
                             in_data[722],
                             in_data[602]};
    
    wire lut_1002_out = lut_1002_table[lut_1002_select];
    
    generate
    if ( USE_REG ) begin : ff_1002
        reg   lut_1002_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1002_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1002_ff <= lut_1002_out;
            end
        end
        
        assign out_data[1002] = lut_1002_ff;
    end
    else begin : no_ff_1002
        assign out_data[1002] = lut_1002_out;
    end
    endgenerate
    
    
    
    // LUT : 1003
    wire [15:0] lut_1003_table = 16'b1110111011101110;
    wire [3:0] lut_1003_select = {
                             in_data[775],
                             in_data[80],
                             in_data[304],
                             in_data[525]};
    
    wire lut_1003_out = lut_1003_table[lut_1003_select];
    
    generate
    if ( USE_REG ) begin : ff_1003
        reg   lut_1003_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1003_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1003_ff <= lut_1003_out;
            end
        end
        
        assign out_data[1003] = lut_1003_ff;
    end
    else begin : no_ff_1003
        assign out_data[1003] = lut_1003_out;
    end
    endgenerate
    
    
    
    // LUT : 1004
    wire [15:0] lut_1004_table = 16'b1101110111011100;
    wire [3:0] lut_1004_select = {
                             in_data[319],
                             in_data[48],
                             in_data[743],
                             in_data[390]};
    
    wire lut_1004_out = lut_1004_table[lut_1004_select];
    
    generate
    if ( USE_REG ) begin : ff_1004
        reg   lut_1004_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1004_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1004_ff <= lut_1004_out;
            end
        end
        
        assign out_data[1004] = lut_1004_ff;
    end
    else begin : no_ff_1004
        assign out_data[1004] = lut_1004_out;
    end
    endgenerate
    
    
    
    // LUT : 1005
    wire [15:0] lut_1005_table = 16'b0101110100000000;
    wire [3:0] lut_1005_select = {
                             in_data[515],
                             in_data[783],
                             in_data[225],
                             in_data[310]};
    
    wire lut_1005_out = lut_1005_table[lut_1005_select];
    
    generate
    if ( USE_REG ) begin : ff_1005
        reg   lut_1005_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1005_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1005_ff <= lut_1005_out;
            end
        end
        
        assign out_data[1005] = lut_1005_ff;
    end
    else begin : no_ff_1005
        assign out_data[1005] = lut_1005_out;
    end
    endgenerate
    
    
    
    // LUT : 1006
    wire [15:0] lut_1006_table = 16'b0000000100000001;
    wire [3:0] lut_1006_select = {
                             in_data[21],
                             in_data[504],
                             in_data[286],
                             in_data[359]};
    
    wire lut_1006_out = lut_1006_table[lut_1006_select];
    
    generate
    if ( USE_REG ) begin : ff_1006
        reg   lut_1006_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1006_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1006_ff <= lut_1006_out;
            end
        end
        
        assign out_data[1006] = lut_1006_ff;
    end
    else begin : no_ff_1006
        assign out_data[1006] = lut_1006_out;
    end
    endgenerate
    
    
    
    // LUT : 1007
    wire [15:0] lut_1007_table = 16'b0010111000111110;
    wire [3:0] lut_1007_select = {
                             in_data[623],
                             in_data[685],
                             in_data[679],
                             in_data[261]};
    
    wire lut_1007_out = lut_1007_table[lut_1007_select];
    
    generate
    if ( USE_REG ) begin : ff_1007
        reg   lut_1007_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1007_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1007_ff <= lut_1007_out;
            end
        end
        
        assign out_data[1007] = lut_1007_ff;
    end
    else begin : no_ff_1007
        assign out_data[1007] = lut_1007_out;
    end
    endgenerate
    
    
    
    // LUT : 1008
    wire [15:0] lut_1008_table = 16'b1111111111001111;
    wire [3:0] lut_1008_select = {
                             in_data[391],
                             in_data[671],
                             in_data[773],
                             in_data[85]};
    
    wire lut_1008_out = lut_1008_table[lut_1008_select];
    
    generate
    if ( USE_REG ) begin : ff_1008
        reg   lut_1008_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1008_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1008_ff <= lut_1008_out;
            end
        end
        
        assign out_data[1008] = lut_1008_ff;
    end
    else begin : no_ff_1008
        assign out_data[1008] = lut_1008_out;
    end
    endgenerate
    
    
    
    // LUT : 1009
    wire [15:0] lut_1009_table = 16'b1111000111110001;
    wire [3:0] lut_1009_select = {
                             in_data[52],
                             in_data[176],
                             in_data[107],
                             in_data[373]};
    
    wire lut_1009_out = lut_1009_table[lut_1009_select];
    
    generate
    if ( USE_REG ) begin : ff_1009
        reg   lut_1009_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1009_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1009_ff <= lut_1009_out;
            end
        end
        
        assign out_data[1009] = lut_1009_ff;
    end
    else begin : no_ff_1009
        assign out_data[1009] = lut_1009_out;
    end
    endgenerate
    
    
    
    // LUT : 1010
    wire [15:0] lut_1010_table = 16'b1111101011111010;
    wire [3:0] lut_1010_select = {
                             in_data[129],
                             in_data[650],
                             in_data[642],
                             in_data[552]};
    
    wire lut_1010_out = lut_1010_table[lut_1010_select];
    
    generate
    if ( USE_REG ) begin : ff_1010
        reg   lut_1010_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1010_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1010_ff <= lut_1010_out;
            end
        end
        
        assign out_data[1010] = lut_1010_ff;
    end
    else begin : no_ff_1010
        assign out_data[1010] = lut_1010_out;
    end
    endgenerate
    
    
    
    // LUT : 1011
    wire [15:0] lut_1011_table = 16'b0000010100000101;
    wire [3:0] lut_1011_select = {
                             in_data[735],
                             in_data[398],
                             in_data[511],
                             in_data[106]};
    
    wire lut_1011_out = lut_1011_table[lut_1011_select];
    
    generate
    if ( USE_REG ) begin : ff_1011
        reg   lut_1011_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1011_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1011_ff <= lut_1011_out;
            end
        end
        
        assign out_data[1011] = lut_1011_ff;
    end
    else begin : no_ff_1011
        assign out_data[1011] = lut_1011_out;
    end
    endgenerate
    
    
    
    // LUT : 1012
    wire [15:0] lut_1012_table = 16'b1111000000110000;
    wire [3:0] lut_1012_select = {
                             in_data[564],
                             in_data[462],
                             in_data[367],
                             in_data[453]};
    
    wire lut_1012_out = lut_1012_table[lut_1012_select];
    
    generate
    if ( USE_REG ) begin : ff_1012
        reg   lut_1012_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1012_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1012_ff <= lut_1012_out;
            end
        end
        
        assign out_data[1012] = lut_1012_ff;
    end
    else begin : no_ff_1012
        assign out_data[1012] = lut_1012_out;
    end
    endgenerate
    
    
    
    // LUT : 1013
    wire [15:0] lut_1013_table = 16'b1011101110101010;
    wire [3:0] lut_1013_select = {
                             in_data[151],
                             in_data[632],
                             in_data[77],
                             in_data[153]};
    
    wire lut_1013_out = lut_1013_table[lut_1013_select];
    
    generate
    if ( USE_REG ) begin : ff_1013
        reg   lut_1013_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1013_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1013_ff <= lut_1013_out;
            end
        end
        
        assign out_data[1013] = lut_1013_ff;
    end
    else begin : no_ff_1013
        assign out_data[1013] = lut_1013_out;
    end
    endgenerate
    
    
    
    // LUT : 1014
    wire [15:0] lut_1014_table = 16'b0011001111001100;
    wire [3:0] lut_1014_select = {
                             in_data[413],
                             in_data[418],
                             in_data[481],
                             in_data[505]};
    
    wire lut_1014_out = lut_1014_table[lut_1014_select];
    
    generate
    if ( USE_REG ) begin : ff_1014
        reg   lut_1014_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1014_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1014_ff <= lut_1014_out;
            end
        end
        
        assign out_data[1014] = lut_1014_ff;
    end
    else begin : no_ff_1014
        assign out_data[1014] = lut_1014_out;
    end
    endgenerate
    
    
    
    // LUT : 1015
    wire [15:0] lut_1015_table = 16'b1111111111110101;
    wire [3:0] lut_1015_select = {
                             in_data[276],
                             in_data[509],
                             in_data[756],
                             in_data[237]};
    
    wire lut_1015_out = lut_1015_table[lut_1015_select];
    
    generate
    if ( USE_REG ) begin : ff_1015
        reg   lut_1015_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1015_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1015_ff <= lut_1015_out;
            end
        end
        
        assign out_data[1015] = lut_1015_ff;
    end
    else begin : no_ff_1015
        assign out_data[1015] = lut_1015_out;
    end
    endgenerate
    
    
    
    // LUT : 1016
    wire [15:0] lut_1016_table = 16'b1111111111111100;
    wire [3:0] lut_1016_select = {
                             in_data[711],
                             in_data[734],
                             in_data[145],
                             in_data[690]};
    
    wire lut_1016_out = lut_1016_table[lut_1016_select];
    
    generate
    if ( USE_REG ) begin : ff_1016
        reg   lut_1016_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1016_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1016_ff <= lut_1016_out;
            end
        end
        
        assign out_data[1016] = lut_1016_ff;
    end
    else begin : no_ff_1016
        assign out_data[1016] = lut_1016_out;
    end
    endgenerate
    
    
    
    // LUT : 1017
    wire [15:0] lut_1017_table = 16'b1011101100110011;
    wire [3:0] lut_1017_select = {
                             in_data[290],
                             in_data[609],
                             in_data[430],
                             in_data[312]};
    
    wire lut_1017_out = lut_1017_table[lut_1017_select];
    
    generate
    if ( USE_REG ) begin : ff_1017
        reg   lut_1017_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1017_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1017_ff <= lut_1017_out;
            end
        end
        
        assign out_data[1017] = lut_1017_ff;
    end
    else begin : no_ff_1017
        assign out_data[1017] = lut_1017_out;
    end
    endgenerate
    
    
    
    // LUT : 1018
    wire [15:0] lut_1018_table = 16'b0011001100000001;
    wire [3:0] lut_1018_select = {
                             in_data[383],
                             in_data[658],
                             in_data[248],
                             in_data[424]};
    
    wire lut_1018_out = lut_1018_table[lut_1018_select];
    
    generate
    if ( USE_REG ) begin : ff_1018
        reg   lut_1018_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1018_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1018_ff <= lut_1018_out;
            end
        end
        
        assign out_data[1018] = lut_1018_ff;
    end
    else begin : no_ff_1018
        assign out_data[1018] = lut_1018_out;
    end
    endgenerate
    
    
    
    // LUT : 1019
    wire [15:0] lut_1019_table = 16'b0000001100101010;
    wire [3:0] lut_1019_select = {
                             in_data[239],
                             in_data[218],
                             in_data[165],
                             in_data[740]};
    
    wire lut_1019_out = lut_1019_table[lut_1019_select];
    
    generate
    if ( USE_REG ) begin : ff_1019
        reg   lut_1019_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1019_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1019_ff <= lut_1019_out;
            end
        end
        
        assign out_data[1019] = lut_1019_ff;
    end
    else begin : no_ff_1019
        assign out_data[1019] = lut_1019_out;
    end
    endgenerate
    
    
    
    // LUT : 1020
    wire [15:0] lut_1020_table = 16'b1111111011111110;
    wire [3:0] lut_1020_select = {
                             in_data[422],
                             in_data[778],
                             in_data[303],
                             in_data[222]};
    
    wire lut_1020_out = lut_1020_table[lut_1020_select];
    
    generate
    if ( USE_REG ) begin : ff_1020
        reg   lut_1020_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1020_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1020_ff <= lut_1020_out;
            end
        end
        
        assign out_data[1020] = lut_1020_ff;
    end
    else begin : no_ff_1020
        assign out_data[1020] = lut_1020_out;
    end
    endgenerate
    
    
    
    // LUT : 1021
    wire [15:0] lut_1021_table = 16'b0011001000110011;
    wire [3:0] lut_1021_select = {
                             in_data[781],
                             in_data[647],
                             in_data[396],
                             in_data[5]};
    
    wire lut_1021_out = lut_1021_table[lut_1021_select];
    
    generate
    if ( USE_REG ) begin : ff_1021
        reg   lut_1021_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1021_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1021_ff <= lut_1021_out;
            end
        end
        
        assign out_data[1021] = lut_1021_ff;
    end
    else begin : no_ff_1021
        assign out_data[1021] = lut_1021_out;
    end
    endgenerate
    
    
    
    // LUT : 1022
    wire [15:0] lut_1022_table = 16'b1010101011111011;
    wire [3:0] lut_1022_select = {
                             in_data[518],
                             in_data[24],
                             in_data[29],
                             in_data[162]};
    
    wire lut_1022_out = lut_1022_table[lut_1022_select];
    
    generate
    if ( USE_REG ) begin : ff_1022
        reg   lut_1022_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1022_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1022_ff <= lut_1022_out;
            end
        end
        
        assign out_data[1022] = lut_1022_ff;
    end
    else begin : no_ff_1022
        assign out_data[1022] = lut_1022_out;
    end
    endgenerate
    
    
    
    // LUT : 1023
    wire [15:0] lut_1023_table = 16'b1111111101010000;
    wire [3:0] lut_1023_select = {
                             in_data[565],
                             in_data[473],
                             in_data[727],
                             in_data[332]};
    
    wire lut_1023_out = lut_1023_table[lut_1023_select];
    
    generate
    if ( USE_REG ) begin : ff_1023
        reg   lut_1023_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1023_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1023_ff <= lut_1023_out;
            end
        end
        
        assign out_data[1023] = lut_1023_ff;
    end
    else begin : no_ff_1023
        assign out_data[1023] = lut_1023_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub1
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [       1023:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        511:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub1_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub1_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub1_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [1023:0]  in_data,
            output wire [511:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1111100000010001;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b1101010111110101;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b1000110100000000;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1100100011001111;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b0000000000010101;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1010101011101111;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b1010111110101111;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1111111111110100;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1111111110100000;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b0001000100010101;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b0000011111111111;
    wire [3:0] lut_10_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b0111001101110011;
    wire [3:0] lut_11_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b1111110011111100;
    wire [3:0] lut_12_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0000000011111111;
    wire [3:0] lut_13_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0010111100100011;
    wire [3:0] lut_14_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1100110011101111;
    wire [3:0] lut_15_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b1010100010110010;
    wire [3:0] lut_16_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b0001011100000101;
    wire [3:0] lut_17_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0000111000011011;
    wire [3:0] lut_18_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b0011001100010001;
    wire [3:0] lut_19_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0101110111011100;
    wire [3:0] lut_20_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b1010101110001111;
    wire [3:0] lut_21_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b1111111100000010;
    wire [3:0] lut_22_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0111010011110100;
    wire [3:0] lut_23_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b0000100010001110;
    wire [3:0] lut_24_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b1111010001010000;
    wire [3:0] lut_25_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b1111000011000000;
    wire [3:0] lut_26_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1111010111010101;
    wire [3:0] lut_27_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b1111010011110101;
    wire [3:0] lut_28_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b0000001100001111;
    wire [3:0] lut_29_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b0001111100001000;
    wire [3:0] lut_30_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1111001001111111;
    wire [3:0] lut_31_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1111000011110000;
    wire [3:0] lut_32_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b1110111100000001;
    wire [3:0] lut_33_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1110000010100000;
    wire [3:0] lut_34_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1101111111001100;
    wire [3:0] lut_35_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b0100010100000000;
    wire [3:0] lut_36_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0000001100010111;
    wire [3:0] lut_37_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b1100101011001100;
    wire [3:0] lut_38_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b1111111100011111;
    wire [3:0] lut_39_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b1111111110001110;
    wire [3:0] lut_40_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b1001000010111011;
    wire [3:0] lut_41_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b1010111110101111;
    wire [3:0] lut_42_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0000000011001100;
    wire [3:0] lut_43_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b0000001111111011;
    wire [3:0] lut_44_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b0101000101011101;
    wire [3:0] lut_45_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b1111001011111111;
    wire [3:0] lut_46_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b0100010011000100;
    wire [3:0] lut_47_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b1010101010101010;
    wire [3:0] lut_48_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b0100000001010000;
    wire [3:0] lut_49_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0101110100011101;
    wire [3:0] lut_50_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b0110000011110111;
    wire [3:0] lut_51_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b0101111100000100;
    wire [3:0] lut_52_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b0011011100100011;
    wire [3:0] lut_53_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b1100110111011101;
    wire [3:0] lut_54_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b0011111100010011;
    wire [3:0] lut_55_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b1000000010110000;
    wire [3:0] lut_56_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b1101111101000101;
    wire [3:0] lut_57_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b0001001100010001;
    wire [3:0] lut_58_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b1100110011001100;
    wire [3:0] lut_59_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b1000000011100000;
    wire [3:0] lut_60_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b0001011100000000;
    wire [3:0] lut_61_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b1100010111001101;
    wire [3:0] lut_62_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b1100111111001111;
    wire [3:0] lut_63_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b1110111111111111;
    wire [3:0] lut_64_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b1010101011100110;
    wire [3:0] lut_65_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b0000111111111111;
    wire [3:0] lut_66_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b1111110111101100;
    wire [3:0] lut_67_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b1111111011110000;
    wire [3:0] lut_68_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b0101111100001111;
    wire [3:0] lut_69_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b0010001000111011;
    wire [3:0] lut_70_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0010111110101111;
    wire [3:0] lut_71_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b0101111101000100;
    wire [3:0] lut_72_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b0000010100000001;
    wire [3:0] lut_73_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0101000001010000;
    wire [3:0] lut_74_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b0000000010101010;
    wire [3:0] lut_75_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0000000001000100;
    wire [3:0] lut_76_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b0101111101011111;
    wire [3:0] lut_77_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b0001010100110001;
    wire [3:0] lut_78_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b0101000001010101;
    wire [3:0] lut_79_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b1111000000001111;
    wire [3:0] lut_80_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b0000000011111011;
    wire [3:0] lut_81_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1111111100001000;
    wire [3:0] lut_82_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b1101110101000101;
    wire [3:0] lut_83_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b0101000000000000;
    wire [3:0] lut_84_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b0000001000111111;
    wire [3:0] lut_85_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b0010111101011111;
    wire [3:0] lut_86_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b1010100010111010;
    wire [3:0] lut_87_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b1010000010000000;
    wire [3:0] lut_88_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b1011001111110001;
    wire [3:0] lut_89_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1110111100001000;
    wire [3:0] lut_90_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b0011000000010000;
    wire [3:0] lut_91_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1111111111001110;
    wire [3:0] lut_92_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0001101000001010;
    wire [3:0] lut_93_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b1101010101010100;
    wire [3:0] lut_94_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b1000001010001010;
    wire [3:0] lut_95_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1111001111110111;
    wire [3:0] lut_96_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b1100000011101100;
    wire [3:0] lut_97_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1111111111110010;
    wire [3:0] lut_98_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b1111000011110101;
    wire [3:0] lut_99_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1010101011001100;
    wire [3:0] lut_100_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b1000110010001100;
    wire [3:0] lut_101_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b0010000011110000;
    wire [3:0] lut_102_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1000110111101111;
    wire [3:0] lut_103_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b0001001000000010;
    wire [3:0] lut_104_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b0000111000001011;
    wire [3:0] lut_105_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b1111010100000000;
    wire [3:0] lut_106_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b0100001001010010;
    wire [3:0] lut_107_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b1101110111000000;
    wire [3:0] lut_108_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b0000111110001111;
    wire [3:0] lut_109_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b1101110111010100;
    wire [3:0] lut_110_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000000001010101;
    wire [3:0] lut_111_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b0111001101111111;
    wire [3:0] lut_112_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b1111111101110011;
    wire [3:0] lut_113_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1111011111111110;
    wire [3:0] lut_114_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0101000110101011;
    wire [3:0] lut_115_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b1111111001001100;
    wire [3:0] lut_116_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b0000111100101011;
    wire [3:0] lut_117_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b0111011100110011;
    wire [3:0] lut_118_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b1111011100000000;
    wire [3:0] lut_119_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b1010011110100111;
    wire [3:0] lut_120_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b0100000111000000;
    wire [3:0] lut_121_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b0101010101110000;
    wire [3:0] lut_122_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b0011111100111111;
    wire [3:0] lut_123_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b1111101011111011;
    wire [3:0] lut_124_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b0111110001010101;
    wire [3:0] lut_125_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b0010010001111111;
    wire [3:0] lut_126_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0000001100011111;
    wire [3:0] lut_127_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b1111111111001111;
    wire [3:0] lut_128_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b0000000000110010;
    wire [3:0] lut_129_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b1111001111110000;
    wire [3:0] lut_130_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b1111000011110001;
    wire [3:0] lut_131_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b1111111100001000;
    wire [3:0] lut_132_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0000000100010111;
    wire [3:0] lut_133_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b1101000011110011;
    wire [3:0] lut_134_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b0111000100010111;
    wire [3:0] lut_135_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b1100100010000000;
    wire [3:0] lut_136_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b0101000000010000;
    wire [3:0] lut_137_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b1111111100100010;
    wire [3:0] lut_138_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b1010101011111111;
    wire [3:0] lut_139_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b0000000000000100;
    wire [3:0] lut_140_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b1111011100010000;
    wire [3:0] lut_141_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b0011000000100000;
    wire [3:0] lut_142_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b1110001010100000;
    wire [3:0] lut_143_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b0111011101110101;
    wire [3:0] lut_144_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1000000010000000;
    wire [3:0] lut_145_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1010000010101010;
    wire [3:0] lut_146_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0000001100111111;
    wire [3:0] lut_147_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b0100000001000100;
    wire [3:0] lut_148_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b1111000011110000;
    wire [3:0] lut_149_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b1100010111111100;
    wire [3:0] lut_150_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b1100000111001111;
    wire [3:0] lut_151_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b0000111100001010;
    wire [3:0] lut_152_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1101111101000000;
    wire [3:0] lut_153_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0111011101110101;
    wire [3:0] lut_154_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b0011001100110010;
    wire [3:0] lut_155_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b0000001100000010;
    wire [3:0] lut_156_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b1111111110101010;
    wire [3:0] lut_157_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b1110000011110000;
    wire [3:0] lut_158_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b0100110101011101;
    wire [3:0] lut_159_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b0000001100111111;
    wire [3:0] lut_160_select = {
                             in_data[643],
                             in_data[642],
                             in_data[641],
                             in_data[640]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b0100110100001100;
    wire [3:0] lut_161_select = {
                             in_data[647],
                             in_data[646],
                             in_data[645],
                             in_data[644]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1110111011111111;
    wire [3:0] lut_162_select = {
                             in_data[651],
                             in_data[650],
                             in_data[649],
                             in_data[648]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b1111111100011111;
    wire [3:0] lut_163_select = {
                             in_data[655],
                             in_data[654],
                             in_data[653],
                             in_data[652]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b1101000111010000;
    wire [3:0] lut_164_select = {
                             in_data[659],
                             in_data[658],
                             in_data[657],
                             in_data[656]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b1010111000000100;
    wire [3:0] lut_165_select = {
                             in_data[663],
                             in_data[662],
                             in_data[661],
                             in_data[660]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b1111000111010100;
    wire [3:0] lut_166_select = {
                             in_data[667],
                             in_data[666],
                             in_data[665],
                             in_data[664]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b0000000001111111;
    wire [3:0] lut_167_select = {
                             in_data[671],
                             in_data[670],
                             in_data[669],
                             in_data[668]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b0101010001000101;
    wire [3:0] lut_168_select = {
                             in_data[675],
                             in_data[674],
                             in_data[673],
                             in_data[672]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b0010101100111011;
    wire [3:0] lut_169_select = {
                             in_data[679],
                             in_data[678],
                             in_data[677],
                             in_data[676]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b1111111111111101;
    wire [3:0] lut_170_select = {
                             in_data[683],
                             in_data[682],
                             in_data[681],
                             in_data[680]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b1010000000000000;
    wire [3:0] lut_171_select = {
                             in_data[687],
                             in_data[686],
                             in_data[685],
                             in_data[684]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b1010001011111111;
    wire [3:0] lut_172_select = {
                             in_data[691],
                             in_data[690],
                             in_data[689],
                             in_data[688]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b1111111111100000;
    wire [3:0] lut_173_select = {
                             in_data[695],
                             in_data[694],
                             in_data[693],
                             in_data[692]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b1011000011110111;
    wire [3:0] lut_174_select = {
                             in_data[699],
                             in_data[698],
                             in_data[697],
                             in_data[696]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1111010111100000;
    wire [3:0] lut_175_select = {
                             in_data[703],
                             in_data[702],
                             in_data[701],
                             in_data[700]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b0000110010001110;
    wire [3:0] lut_176_select = {
                             in_data[707],
                             in_data[706],
                             in_data[705],
                             in_data[704]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b0000111000111111;
    wire [3:0] lut_177_select = {
                             in_data[711],
                             in_data[710],
                             in_data[709],
                             in_data[708]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b1000111110001111;
    wire [3:0] lut_178_select = {
                             in_data[715],
                             in_data[714],
                             in_data[713],
                             in_data[712]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b0011001000001011;
    wire [3:0] lut_179_select = {
                             in_data[719],
                             in_data[718],
                             in_data[717],
                             in_data[716]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b1111111111110000;
    wire [3:0] lut_180_select = {
                             in_data[723],
                             in_data[722],
                             in_data[721],
                             in_data[720]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b1101111101011101;
    wire [3:0] lut_181_select = {
                             in_data[727],
                             in_data[726],
                             in_data[725],
                             in_data[724]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b1010101110000011;
    wire [3:0] lut_182_select = {
                             in_data[731],
                             in_data[730],
                             in_data[729],
                             in_data[728]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b1111001111110011;
    wire [3:0] lut_183_select = {
                             in_data[735],
                             in_data[734],
                             in_data[733],
                             in_data[732]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b1111110011000000;
    wire [3:0] lut_184_select = {
                             in_data[739],
                             in_data[738],
                             in_data[737],
                             in_data[736]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b0000000001111111;
    wire [3:0] lut_185_select = {
                             in_data[743],
                             in_data[742],
                             in_data[741],
                             in_data[740]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b0101010101010111;
    wire [3:0] lut_186_select = {
                             in_data[747],
                             in_data[746],
                             in_data[745],
                             in_data[744]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b0000101000001111;
    wire [3:0] lut_187_select = {
                             in_data[751],
                             in_data[750],
                             in_data[749],
                             in_data[748]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b0000000001011101;
    wire [3:0] lut_188_select = {
                             in_data[755],
                             in_data[754],
                             in_data[753],
                             in_data[752]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b0010101100000000;
    wire [3:0] lut_189_select = {
                             in_data[759],
                             in_data[758],
                             in_data[757],
                             in_data[756]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b1111011111110111;
    wire [3:0] lut_190_select = {
                             in_data[763],
                             in_data[762],
                             in_data[761],
                             in_data[760]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b1111110011010101;
    wire [3:0] lut_191_select = {
                             in_data[767],
                             in_data[766],
                             in_data[765],
                             in_data[764]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b1010111111001111;
    wire [3:0] lut_192_select = {
                             in_data[771],
                             in_data[770],
                             in_data[769],
                             in_data[768]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b0111001101110011;
    wire [3:0] lut_193_select = {
                             in_data[775],
                             in_data[774],
                             in_data[773],
                             in_data[772]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0101010101010101;
    wire [3:0] lut_194_select = {
                             in_data[779],
                             in_data[778],
                             in_data[777],
                             in_data[776]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b0100110000001111;
    wire [3:0] lut_195_select = {
                             in_data[783],
                             in_data[782],
                             in_data[781],
                             in_data[780]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b0101100001001000;
    wire [3:0] lut_196_select = {
                             in_data[787],
                             in_data[786],
                             in_data[785],
                             in_data[784]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b1000110000000000;
    wire [3:0] lut_197_select = {
                             in_data[791],
                             in_data[790],
                             in_data[789],
                             in_data[788]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b1010111000000000;
    wire [3:0] lut_198_select = {
                             in_data[795],
                             in_data[794],
                             in_data[793],
                             in_data[792]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b1111010111110111;
    wire [3:0] lut_199_select = {
                             in_data[799],
                             in_data[798],
                             in_data[797],
                             in_data[796]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b0011101100111011;
    wire [3:0] lut_200_select = {
                             in_data[803],
                             in_data[802],
                             in_data[801],
                             in_data[800]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b1101111111011100;
    wire [3:0] lut_201_select = {
                             in_data[807],
                             in_data[806],
                             in_data[805],
                             in_data[804]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b1000110010001110;
    wire [3:0] lut_202_select = {
                             in_data[811],
                             in_data[810],
                             in_data[809],
                             in_data[808]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b0000001110000011;
    wire [3:0] lut_203_select = {
                             in_data[815],
                             in_data[814],
                             in_data[813],
                             in_data[812]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b1101000011111101;
    wire [3:0] lut_204_select = {
                             in_data[819],
                             in_data[818],
                             in_data[817],
                             in_data[816]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b1111000011110000;
    wire [3:0] lut_205_select = {
                             in_data[823],
                             in_data[822],
                             in_data[821],
                             in_data[820]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b1010101010101010;
    wire [3:0] lut_206_select = {
                             in_data[827],
                             in_data[826],
                             in_data[825],
                             in_data[824]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b0000011100000001;
    wire [3:0] lut_207_select = {
                             in_data[831],
                             in_data[830],
                             in_data[829],
                             in_data[828]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1111111101000101;
    wire [3:0] lut_208_select = {
                             in_data[835],
                             in_data[834],
                             in_data[833],
                             in_data[832]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b0001001100000000;
    wire [3:0] lut_209_select = {
                             in_data[839],
                             in_data[838],
                             in_data[837],
                             in_data[836]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b1010111010110011;
    wire [3:0] lut_210_select = {
                             in_data[843],
                             in_data[842],
                             in_data[841],
                             in_data[840]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b1101110100000000;
    wire [3:0] lut_211_select = {
                             in_data[847],
                             in_data[846],
                             in_data[845],
                             in_data[844]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b0100000000010001;
    wire [3:0] lut_212_select = {
                             in_data[851],
                             in_data[850],
                             in_data[849],
                             in_data[848]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b0101010001000101;
    wire [3:0] lut_213_select = {
                             in_data[855],
                             in_data[854],
                             in_data[853],
                             in_data[852]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1000001011001111;
    wire [3:0] lut_214_select = {
                             in_data[859],
                             in_data[858],
                             in_data[857],
                             in_data[856]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b1111111111111010;
    wire [3:0] lut_215_select = {
                             in_data[863],
                             in_data[862],
                             in_data[861],
                             in_data[860]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b0011011101000100;
    wire [3:0] lut_216_select = {
                             in_data[867],
                             in_data[866],
                             in_data[865],
                             in_data[864]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b0111011111110000;
    wire [3:0] lut_217_select = {
                             in_data[871],
                             in_data[870],
                             in_data[869],
                             in_data[868]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b1000000010100010;
    wire [3:0] lut_218_select = {
                             in_data[875],
                             in_data[874],
                             in_data[873],
                             in_data[872]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b1111111111011111;
    wire [3:0] lut_219_select = {
                             in_data[879],
                             in_data[878],
                             in_data[877],
                             in_data[876]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b1101010011110101;
    wire [3:0] lut_220_select = {
                             in_data[883],
                             in_data[882],
                             in_data[881],
                             in_data[880]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b0010011000111110;
    wire [3:0] lut_221_select = {
                             in_data[887],
                             in_data[886],
                             in_data[885],
                             in_data[884]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b0101110001010000;
    wire [3:0] lut_222_select = {
                             in_data[891],
                             in_data[890],
                             in_data[889],
                             in_data[888]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1111111111011100;
    wire [3:0] lut_223_select = {
                             in_data[895],
                             in_data[894],
                             in_data[893],
                             in_data[892]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b0111000011111111;
    wire [3:0] lut_224_select = {
                             in_data[899],
                             in_data[898],
                             in_data[897],
                             in_data[896]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b1111101011110010;
    wire [3:0] lut_225_select = {
                             in_data[903],
                             in_data[902],
                             in_data[901],
                             in_data[900]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1111010111110100;
    wire [3:0] lut_226_select = {
                             in_data[907],
                             in_data[906],
                             in_data[905],
                             in_data[904]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b1000100011001100;
    wire [3:0] lut_227_select = {
                             in_data[911],
                             in_data[910],
                             in_data[909],
                             in_data[908]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b1010110000001100;
    wire [3:0] lut_228_select = {
                             in_data[915],
                             in_data[914],
                             in_data[913],
                             in_data[912]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b1111111111001111;
    wire [3:0] lut_229_select = {
                             in_data[919],
                             in_data[918],
                             in_data[917],
                             in_data[916]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b0000000011001100;
    wire [3:0] lut_230_select = {
                             in_data[923],
                             in_data[922],
                             in_data[921],
                             in_data[920]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b0111001100110010;
    wire [3:0] lut_231_select = {
                             in_data[927],
                             in_data[926],
                             in_data[925],
                             in_data[924]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b0111001100110011;
    wire [3:0] lut_232_select = {
                             in_data[931],
                             in_data[930],
                             in_data[929],
                             in_data[928]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b1000110011001101;
    wire [3:0] lut_233_select = {
                             in_data[935],
                             in_data[934],
                             in_data[933],
                             in_data[932]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b1111111011101010;
    wire [3:0] lut_234_select = {
                             in_data[939],
                             in_data[938],
                             in_data[937],
                             in_data[936]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b0100010011010100;
    wire [3:0] lut_235_select = {
                             in_data[943],
                             in_data[942],
                             in_data[941],
                             in_data[940]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b1011001010111111;
    wire [3:0] lut_236_select = {
                             in_data[947],
                             in_data[946],
                             in_data[945],
                             in_data[944]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b0000011100001111;
    wire [3:0] lut_237_select = {
                             in_data[951],
                             in_data[950],
                             in_data[949],
                             in_data[948]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b0100010011100100;
    wire [3:0] lut_238_select = {
                             in_data[955],
                             in_data[954],
                             in_data[953],
                             in_data[952]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0000010000001111;
    wire [3:0] lut_239_select = {
                             in_data[959],
                             in_data[958],
                             in_data[957],
                             in_data[956]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b0101010011010000;
    wire [3:0] lut_240_select = {
                             in_data[963],
                             in_data[962],
                             in_data[961],
                             in_data[960]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b1110111011111110;
    wire [3:0] lut_241_select = {
                             in_data[967],
                             in_data[966],
                             in_data[965],
                             in_data[964]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b0101000001010000;
    wire [3:0] lut_242_select = {
                             in_data[971],
                             in_data[970],
                             in_data[969],
                             in_data[968]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b0000111011111111;
    wire [3:0] lut_243_select = {
                             in_data[975],
                             in_data[974],
                             in_data[973],
                             in_data[972]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b1010101011111111;
    wire [3:0] lut_244_select = {
                             in_data[979],
                             in_data[978],
                             in_data[977],
                             in_data[976]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b0101011100010000;
    wire [3:0] lut_245_select = {
                             in_data[983],
                             in_data[982],
                             in_data[981],
                             in_data[980]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b0000110000000011;
    wire [3:0] lut_246_select = {
                             in_data[987],
                             in_data[986],
                             in_data[985],
                             in_data[984]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b0000000100010101;
    wire [3:0] lut_247_select = {
                             in_data[991],
                             in_data[990],
                             in_data[989],
                             in_data[988]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b0000100010001111;
    wire [3:0] lut_248_select = {
                             in_data[995],
                             in_data[994],
                             in_data[993],
                             in_data[992]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b0001000000000000;
    wire [3:0] lut_249_select = {
                             in_data[999],
                             in_data[998],
                             in_data[997],
                             in_data[996]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b0000001100101011;
    wire [3:0] lut_250_select = {
                             in_data[1003],
                             in_data[1002],
                             in_data[1001],
                             in_data[1000]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b0000000011110000;
    wire [3:0] lut_251_select = {
                             in_data[1007],
                             in_data[1006],
                             in_data[1005],
                             in_data[1004]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b0001000101010101;
    wire [3:0] lut_252_select = {
                             in_data[1011],
                             in_data[1010],
                             in_data[1009],
                             in_data[1008]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b1011101110101000;
    wire [3:0] lut_253_select = {
                             in_data[1015],
                             in_data[1014],
                             in_data[1013],
                             in_data[1012]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b1110111110001000;
    wire [3:0] lut_254_select = {
                             in_data[1019],
                             in_data[1018],
                             in_data[1017],
                             in_data[1016]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b1100110100000100;
    wire [3:0] lut_255_select = {
                             in_data[1023],
                             in_data[1022],
                             in_data[1021],
                             in_data[1020]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b0100010101011111;
    wire [3:0] lut_256_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b0010001000001111;
    wire [3:0] lut_257_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b1101110011111110;
    wire [3:0] lut_258_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b0111001100110001;
    wire [3:0] lut_259_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b1111000010110000;
    wire [3:0] lut_260_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b0001000100110001;
    wire [3:0] lut_261_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b0000110100000101;
    wire [3:0] lut_262_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b0000000011110001;
    wire [3:0] lut_263_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b1111111111001010;
    wire [3:0] lut_264_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b1111110011000000;
    wire [3:0] lut_265_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1111000000000101;
    wire [3:0] lut_266_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b1100010011111100;
    wire [3:0] lut_267_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1000100010001110;
    wire [3:0] lut_268_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0111000011110000;
    wire [3:0] lut_269_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b0001111100011111;
    wire [3:0] lut_270_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b0000110010001110;
    wire [3:0] lut_271_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b0011101100110011;
    wire [3:0] lut_272_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b0111111100000101;
    wire [3:0] lut_273_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b1111111111100100;
    wire [3:0] lut_274_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b0101000101010001;
    wire [3:0] lut_275_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b0000101011110000;
    wire [3:0] lut_276_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b0111010100000000;
    wire [3:0] lut_277_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b1111111110110011;
    wire [3:0] lut_278_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b0011111100111111;
    wire [3:0] lut_279_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b1111001101110001;
    wire [3:0] lut_280_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b0111010100010000;
    wire [3:0] lut_281_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b1111000011000000;
    wire [3:0] lut_282_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b1101001100000010;
    wire [3:0] lut_283_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b0000111000001110;
    wire [3:0] lut_284_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b0000110100001111;
    wire [3:0] lut_285_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b0111111110001000;
    wire [3:0] lut_286_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b0010000000100011;
    wire [3:0] lut_287_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b0111011101010001;
    wire [3:0] lut_288_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b0111111100010011;
    wire [3:0] lut_289_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b0001000100011111;
    wire [3:0] lut_290_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b0111000011111010;
    wire [3:0] lut_291_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b1111010100000000;
    wire [3:0] lut_292_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b0011101100111111;
    wire [3:0] lut_293_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1011001100000010;
    wire [3:0] lut_294_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b0000010101001101;
    wire [3:0] lut_295_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b1110111011101110;
    wire [3:0] lut_296_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b0100111101000000;
    wire [3:0] lut_297_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b1011111100101111;
    wire [3:0] lut_298_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b1000000011001100;
    wire [3:0] lut_299_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b0010001011110010;
    wire [3:0] lut_300_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b0100010111111111;
    wire [3:0] lut_301_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b0000010001011111;
    wire [3:0] lut_302_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b1011101100101011;
    wire [3:0] lut_303_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b0100010101000101;
    wire [3:0] lut_304_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b0001000001010000;
    wire [3:0] lut_305_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b0101010101010101;
    wire [3:0] lut_306_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b1010000011111100;
    wire [3:0] lut_307_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b1111001011100010;
    wire [3:0] lut_308_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b0111000000110010;
    wire [3:0] lut_309_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b0011001000100010;
    wire [3:0] lut_310_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b0100000001110000;
    wire [3:0] lut_311_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1000000010000000;
    wire [3:0] lut_312_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b1101110101010101;
    wire [3:0] lut_313_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b0101010100010101;
    wire [3:0] lut_314_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b1101000100110000;
    wire [3:0] lut_315_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b1011001100110011;
    wire [3:0] lut_316_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b1110111011111111;
    wire [3:0] lut_317_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0000000011110101;
    wire [3:0] lut_318_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b1011001010110000;
    wire [3:0] lut_319_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b1110111111111111;
    wire [3:0] lut_320_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0001000100010001;
    wire [3:0] lut_321_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b1100110011111111;
    wire [3:0] lut_322_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b0011111100010101;
    wire [3:0] lut_323_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b0000010100000101;
    wire [3:0] lut_324_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b1010000000100000;
    wire [3:0] lut_325_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b0000010011010101;
    wire [3:0] lut_326_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b0000000010101010;
    wire [3:0] lut_327_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b0000001000000000;
    wire [3:0] lut_328_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b0000110101001101;
    wire [3:0] lut_329_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b0100000011001100;
    wire [3:0] lut_330_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b1000111100001111;
    wire [3:0] lut_331_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b0001011101110111;
    wire [3:0] lut_332_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b1010000010100000;
    wire [3:0] lut_333_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b0000010100010001;
    wire [3:0] lut_334_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0100010001000100;
    wire [3:0] lut_335_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b0011111100110000;
    wire [3:0] lut_336_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b0000000000000001;
    wire [3:0] lut_337_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b1111011100000000;
    wire [3:0] lut_338_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b1111010101010000;
    wire [3:0] lut_339_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b1010111110111111;
    wire [3:0] lut_340_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b0111000100010000;
    wire [3:0] lut_341_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b1101100000000000;
    wire [3:0] lut_342_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b1000100010101010;
    wire [3:0] lut_343_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1010100000000000;
    wire [3:0] lut_344_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b1111111101010101;
    wire [3:0] lut_345_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b1101000000000000;
    wire [3:0] lut_346_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b0011000000000000;
    wire [3:0] lut_347_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0000000000110001;
    wire [3:0] lut_348_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b1000100010001000;
    wire [3:0] lut_349_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b0101010111010101;
    wire [3:0] lut_350_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b0011000101110001;
    wire [3:0] lut_351_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b1111111110110011;
    wire [3:0] lut_352_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b0000000010001000;
    wire [3:0] lut_353_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b0000010001000101;
    wire [3:0] lut_354_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b0000111110001100;
    wire [3:0] lut_355_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b1010101001001100;
    wire [3:0] lut_356_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b0011111111111101;
    wire [3:0] lut_357_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b1010111100001111;
    wire [3:0] lut_358_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b1100111111001101;
    wire [3:0] lut_359_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b0000011011101110;
    wire [3:0] lut_360_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b0111010100100000;
    wire [3:0] lut_361_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b1111010100000000;
    wire [3:0] lut_362_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b1010000011101110;
    wire [3:0] lut_363_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b1101010111001000;
    wire [3:0] lut_364_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b0000111111001111;
    wire [3:0] lut_365_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b1101110111010000;
    wire [3:0] lut_366_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b1011000110001000;
    wire [3:0] lut_367_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b1000110010001000;
    wire [3:0] lut_368_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b1000000011001000;
    wire [3:0] lut_369_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b1111111111110110;
    wire [3:0] lut_370_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b0000010110111111;
    wire [3:0] lut_371_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b1111011001001100;
    wire [3:0] lut_372_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b1111110011111000;
    wire [3:0] lut_373_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b1110100011001100;
    wire [3:0] lut_374_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b1100111000001100;
    wire [3:0] lut_375_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b1110011111000111;
    wire [3:0] lut_376_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b1111011100000001;
    wire [3:0] lut_377_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b1010101010101111;
    wire [3:0] lut_378_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1101110111010001;
    wire [3:0] lut_379_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b0100010001000100;
    wire [3:0] lut_380_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b0100110101001101;
    wire [3:0] lut_381_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b0101011101110111;
    wire [3:0] lut_382_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b1101110101010101;
    wire [3:0] lut_383_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0111111111001111;
    wire [3:0] lut_384_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b1101011101000101;
    wire [3:0] lut_385_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b1111101111110011;
    wire [3:0] lut_386_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b1111011100010001;
    wire [3:0] lut_387_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b1000101110001110;
    wire [3:0] lut_388_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b1111111101000000;
    wire [3:0] lut_389_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b0101010101000101;
    wire [3:0] lut_390_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b0011000100010111;
    wire [3:0] lut_391_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b0011000100111011;
    wire [3:0] lut_392_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b0011000100010000;
    wire [3:0] lut_393_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b0010101000001010;
    wire [3:0] lut_394_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b1000110100000000;
    wire [3:0] lut_395_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b0000100000001010;
    wire [3:0] lut_396_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b0000111110001111;
    wire [3:0] lut_397_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b1111001001000000;
    wire [3:0] lut_398_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b0000000000111011;
    wire [3:0] lut_399_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b0111011111110111;
    wire [3:0] lut_400_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b0001111100011111;
    wire [3:0] lut_401_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b0000000010101010;
    wire [3:0] lut_402_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b0100110000000000;
    wire [3:0] lut_403_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b1011101110110010;
    wire [3:0] lut_404_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b0100100001011000;
    wire [3:0] lut_405_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0000110100001111;
    wire [3:0] lut_406_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b1100101111001111;
    wire [3:0] lut_407_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b0000001100010011;
    wire [3:0] lut_408_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b0101000001010100;
    wire [3:0] lut_409_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b1111111111110000;
    wire [3:0] lut_410_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b0101010101010101;
    wire [3:0] lut_411_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b0000111000111111;
    wire [3:0] lut_412_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b0001000011110101;
    wire [3:0] lut_413_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0101001101000001;
    wire [3:0] lut_414_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b1011111100001101;
    wire [3:0] lut_415_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b1011001111111011;
    wire [3:0] lut_416_select = {
                             in_data[643],
                             in_data[642],
                             in_data[641],
                             in_data[640]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b1010000011110010;
    wire [3:0] lut_417_select = {
                             in_data[647],
                             in_data[646],
                             in_data[645],
                             in_data[644]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b1110111011111111;
    wire [3:0] lut_418_select = {
                             in_data[651],
                             in_data[650],
                             in_data[649],
                             in_data[648]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b1111111110111111;
    wire [3:0] lut_419_select = {
                             in_data[655],
                             in_data[654],
                             in_data[653],
                             in_data[652]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b1010101000010000;
    wire [3:0] lut_420_select = {
                             in_data[659],
                             in_data[658],
                             in_data[657],
                             in_data[656]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b0111001111111111;
    wire [3:0] lut_421_select = {
                             in_data[663],
                             in_data[662],
                             in_data[661],
                             in_data[660]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b1101010011111100;
    wire [3:0] lut_422_select = {
                             in_data[667],
                             in_data[666],
                             in_data[665],
                             in_data[664]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b0000000111111111;
    wire [3:0] lut_423_select = {
                             in_data[671],
                             in_data[670],
                             in_data[669],
                             in_data[668]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b0001000011010000;
    wire [3:0] lut_424_select = {
                             in_data[675],
                             in_data[674],
                             in_data[673],
                             in_data[672]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b0000000010100010;
    wire [3:0] lut_425_select = {
                             in_data[679],
                             in_data[678],
                             in_data[677],
                             in_data[676]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b0000000000100010;
    wire [3:0] lut_426_select = {
                             in_data[683],
                             in_data[682],
                             in_data[681],
                             in_data[680]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b0101111111111011;
    wire [3:0] lut_427_select = {
                             in_data[687],
                             in_data[686],
                             in_data[685],
                             in_data[684]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b0000000000000011;
    wire [3:0] lut_428_select = {
                             in_data[691],
                             in_data[690],
                             in_data[689],
                             in_data[688]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b0000110111111111;
    wire [3:0] lut_429_select = {
                             in_data[695],
                             in_data[694],
                             in_data[693],
                             in_data[692]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b0011001111110111;
    wire [3:0] lut_430_select = {
                             in_data[699],
                             in_data[698],
                             in_data[697],
                             in_data[696]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b0010101100011111;
    wire [3:0] lut_431_select = {
                             in_data[703],
                             in_data[702],
                             in_data[701],
                             in_data[700]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b0000100000001111;
    wire [3:0] lut_432_select = {
                             in_data[707],
                             in_data[706],
                             in_data[705],
                             in_data[704]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b1100000000000000;
    wire [3:0] lut_433_select = {
                             in_data[711],
                             in_data[710],
                             in_data[709],
                             in_data[708]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b1000111110001101;
    wire [3:0] lut_434_select = {
                             in_data[715],
                             in_data[714],
                             in_data[713],
                             in_data[712]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b0001001010001010;
    wire [3:0] lut_435_select = {
                             in_data[719],
                             in_data[718],
                             in_data[717],
                             in_data[716]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b1101000011110000;
    wire [3:0] lut_436_select = {
                             in_data[723],
                             in_data[722],
                             in_data[721],
                             in_data[720]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b0001010100010101;
    wire [3:0] lut_437_select = {
                             in_data[727],
                             in_data[726],
                             in_data[725],
                             in_data[724]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b0101100000001000;
    wire [3:0] lut_438_select = {
                             in_data[731],
                             in_data[730],
                             in_data[729],
                             in_data[728]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b0101010101011101;
    wire [3:0] lut_439_select = {
                             in_data[735],
                             in_data[734],
                             in_data[733],
                             in_data[732]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b0011001110111111;
    wire [3:0] lut_440_select = {
                             in_data[739],
                             in_data[738],
                             in_data[737],
                             in_data[736]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b1000111010101010;
    wire [3:0] lut_441_select = {
                             in_data[743],
                             in_data[742],
                             in_data[741],
                             in_data[740]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b1010101010000000;
    wire [3:0] lut_442_select = {
                             in_data[747],
                             in_data[746],
                             in_data[745],
                             in_data[744]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1111000001010000;
    wire [3:0] lut_443_select = {
                             in_data[751],
                             in_data[750],
                             in_data[749],
                             in_data[748]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b0100111101001101;
    wire [3:0] lut_444_select = {
                             in_data[755],
                             in_data[754],
                             in_data[753],
                             in_data[752]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b1110101011001000;
    wire [3:0] lut_445_select = {
                             in_data[759],
                             in_data[758],
                             in_data[757],
                             in_data[756]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b1010101110111011;
    wire [3:0] lut_446_select = {
                             in_data[763],
                             in_data[762],
                             in_data[761],
                             in_data[760]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b0101010110111011;
    wire [3:0] lut_447_select = {
                             in_data[767],
                             in_data[766],
                             in_data[765],
                             in_data[764]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b0001000000110001;
    wire [3:0] lut_448_select = {
                             in_data[771],
                             in_data[770],
                             in_data[769],
                             in_data[768]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b0000110100001101;
    wire [3:0] lut_449_select = {
                             in_data[775],
                             in_data[774],
                             in_data[773],
                             in_data[772]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b1110100011101000;
    wire [3:0] lut_450_select = {
                             in_data[779],
                             in_data[778],
                             in_data[777],
                             in_data[776]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b1011101111111111;
    wire [3:0] lut_451_select = {
                             in_data[783],
                             in_data[782],
                             in_data[781],
                             in_data[780]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b0101100001001000;
    wire [3:0] lut_452_select = {
                             in_data[787],
                             in_data[786],
                             in_data[785],
                             in_data[784]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b1000110000000000;
    wire [3:0] lut_453_select = {
                             in_data[791],
                             in_data[790],
                             in_data[789],
                             in_data[788]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0101000111111111;
    wire [3:0] lut_454_select = {
                             in_data[795],
                             in_data[794],
                             in_data[793],
                             in_data[792]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b0000101000000000;
    wire [3:0] lut_455_select = {
                             in_data[799],
                             in_data[798],
                             in_data[797],
                             in_data[796]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b1011111100101011;
    wire [3:0] lut_456_select = {
                             in_data[803],
                             in_data[802],
                             in_data[801],
                             in_data[800]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b0100110101011101;
    wire [3:0] lut_457_select = {
                             in_data[807],
                             in_data[806],
                             in_data[805],
                             in_data[804]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b1100000010000000;
    wire [3:0] lut_458_select = {
                             in_data[811],
                             in_data[810],
                             in_data[809],
                             in_data[808]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b1100110111001111;
    wire [3:0] lut_459_select = {
                             in_data[815],
                             in_data[814],
                             in_data[813],
                             in_data[812]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b1100110100011111;
    wire [3:0] lut_460_select = {
                             in_data[819],
                             in_data[818],
                             in_data[817],
                             in_data[816]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b1101000011011100;
    wire [3:0] lut_461_select = {
                             in_data[823],
                             in_data[822],
                             in_data[821],
                             in_data[820]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b1000110010001100;
    wire [3:0] lut_462_select = {
                             in_data[827],
                             in_data[826],
                             in_data[825],
                             in_data[824]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b0001000011111011;
    wire [3:0] lut_463_select = {
                             in_data[831],
                             in_data[830],
                             in_data[829],
                             in_data[828]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b0000111111001111;
    wire [3:0] lut_464_select = {
                             in_data[835],
                             in_data[834],
                             in_data[833],
                             in_data[832]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b0011001111110011;
    wire [3:0] lut_465_select = {
                             in_data[839],
                             in_data[838],
                             in_data[837],
                             in_data[836]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b1000111110100001;
    wire [3:0] lut_466_select = {
                             in_data[843],
                             in_data[842],
                             in_data[841],
                             in_data[840]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1100110011000000;
    wire [3:0] lut_467_select = {
                             in_data[847],
                             in_data[846],
                             in_data[845],
                             in_data[844]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b0001011101111111;
    wire [3:0] lut_468_select = {
                             in_data[851],
                             in_data[850],
                             in_data[849],
                             in_data[848]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b0000111100001111;
    wire [3:0] lut_469_select = {
                             in_data[855],
                             in_data[854],
                             in_data[853],
                             in_data[852]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b1011100010111000;
    wire [3:0] lut_470_select = {
                             in_data[859],
                             in_data[858],
                             in_data[857],
                             in_data[856]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b0010000011110000;
    wire [3:0] lut_471_select = {
                             in_data[863],
                             in_data[862],
                             in_data[861],
                             in_data[860]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b1100111011001100;
    wire [3:0] lut_472_select = {
                             in_data[867],
                             in_data[866],
                             in_data[865],
                             in_data[864]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b0000110000001111;
    wire [3:0] lut_473_select = {
                             in_data[871],
                             in_data[870],
                             in_data[869],
                             in_data[868]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b0101110101000101;
    wire [3:0] lut_474_select = {
                             in_data[875],
                             in_data[874],
                             in_data[873],
                             in_data[872]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b0000000000110000;
    wire [3:0] lut_475_select = {
                             in_data[879],
                             in_data[878],
                             in_data[877],
                             in_data[876]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b0010001000101010;
    wire [3:0] lut_476_select = {
                             in_data[883],
                             in_data[882],
                             in_data[881],
                             in_data[880]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b1101000011000000;
    wire [3:0] lut_477_select = {
                             in_data[887],
                             in_data[886],
                             in_data[885],
                             in_data[884]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b0010101100101011;
    wire [3:0] lut_478_select = {
                             in_data[891],
                             in_data[890],
                             in_data[889],
                             in_data[888]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b1111111100001010;
    wire [3:0] lut_479_select = {
                             in_data[895],
                             in_data[894],
                             in_data[893],
                             in_data[892]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b1111001111111111;
    wire [3:0] lut_480_select = {
                             in_data[899],
                             in_data[898],
                             in_data[897],
                             in_data[896]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b0000010100001101;
    wire [3:0] lut_481_select = {
                             in_data[903],
                             in_data[902],
                             in_data[901],
                             in_data[900]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b0000100010001111;
    wire [3:0] lut_482_select = {
                             in_data[907],
                             in_data[906],
                             in_data[905],
                             in_data[904]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b1000100011001100;
    wire [3:0] lut_483_select = {
                             in_data[911],
                             in_data[910],
                             in_data[909],
                             in_data[908]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b0011001101110011;
    wire [3:0] lut_484_select = {
                             in_data[915],
                             in_data[914],
                             in_data[913],
                             in_data[912]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b0000000001110011;
    wire [3:0] lut_485_select = {
                             in_data[919],
                             in_data[918],
                             in_data[917],
                             in_data[916]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b0101010111011101;
    wire [3:0] lut_486_select = {
                             in_data[923],
                             in_data[922],
                             in_data[921],
                             in_data[920]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b1000000000000000;
    wire [3:0] lut_487_select = {
                             in_data[927],
                             in_data[926],
                             in_data[925],
                             in_data[924]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1111010111110101;
    wire [3:0] lut_488_select = {
                             in_data[931],
                             in_data[930],
                             in_data[929],
                             in_data[928]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b0111101000001010;
    wire [3:0] lut_489_select = {
                             in_data[935],
                             in_data[934],
                             in_data[933],
                             in_data[932]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b1110111011101110;
    wire [3:0] lut_490_select = {
                             in_data[939],
                             in_data[938],
                             in_data[937],
                             in_data[936]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b1010111110001110;
    wire [3:0] lut_491_select = {
                             in_data[943],
                             in_data[942],
                             in_data[941],
                             in_data[940]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b1000000011001100;
    wire [3:0] lut_492_select = {
                             in_data[947],
                             in_data[946],
                             in_data[945],
                             in_data[944]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b1100110111001111;
    wire [3:0] lut_493_select = {
                             in_data[951],
                             in_data[950],
                             in_data[949],
                             in_data[948]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b1111111011101100;
    wire [3:0] lut_494_select = {
                             in_data[955],
                             in_data[954],
                             in_data[953],
                             in_data[952]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b0000010000001111;
    wire [3:0] lut_495_select = {
                             in_data[959],
                             in_data[958],
                             in_data[957],
                             in_data[956]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b1101110111001100;
    wire [3:0] lut_496_select = {
                             in_data[963],
                             in_data[962],
                             in_data[961],
                             in_data[960]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b1010111111101110;
    wire [3:0] lut_497_select = {
                             in_data[967],
                             in_data[966],
                             in_data[965],
                             in_data[964]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b1010111111101111;
    wire [3:0] lut_498_select = {
                             in_data[971],
                             in_data[970],
                             in_data[969],
                             in_data[968]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b0000101011111010;
    wire [3:0] lut_499_select = {
                             in_data[975],
                             in_data[974],
                             in_data[973],
                             in_data[972]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b0111000100000000;
    wire [3:0] lut_500_select = {
                             in_data[979],
                             in_data[978],
                             in_data[977],
                             in_data[976]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b0001011100000000;
    wire [3:0] lut_501_select = {
                             in_data[983],
                             in_data[982],
                             in_data[981],
                             in_data[980]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b0000100000001000;
    wire [3:0] lut_502_select = {
                             in_data[987],
                             in_data[986],
                             in_data[985],
                             in_data[984]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b1111111011101000;
    wire [3:0] lut_503_select = {
                             in_data[991],
                             in_data[990],
                             in_data[989],
                             in_data[988]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b1111111111110101;
    wire [3:0] lut_504_select = {
                             in_data[995],
                             in_data[994],
                             in_data[993],
                             in_data[992]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b0011000011110000;
    wire [3:0] lut_505_select = {
                             in_data[999],
                             in_data[998],
                             in_data[997],
                             in_data[996]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b0001000011110000;
    wire [3:0] lut_506_select = {
                             in_data[1003],
                             in_data[1002],
                             in_data[1001],
                             in_data[1000]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b1100110011001100;
    wire [3:0] lut_507_select = {
                             in_data[1007],
                             in_data[1006],
                             in_data[1005],
                             in_data[1004]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b1111110010110010;
    wire [3:0] lut_508_select = {
                             in_data[1011],
                             in_data[1010],
                             in_data[1009],
                             in_data[1008]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b0101000101010111;
    wire [3:0] lut_509_select = {
                             in_data[1015],
                             in_data[1014],
                             in_data[1013],
                             in_data[1012]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b0000010101110111;
    wire [3:0] lut_510_select = {
                             in_data[1019],
                             in_data[1018],
                             in_data[1017],
                             in_data[1016]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0000000000111111;
    wire [3:0] lut_511_select = {
                             in_data[1023],
                             in_data[1022],
                             in_data[1021],
                             in_data[1020]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub2
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        511:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        639:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub2_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub2_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub2_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [511:0]  in_data,
            output wire [639:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1111001111110010;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b0111010111110111;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b1000000011111011;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b0111111101110111;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b0010001100111011;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b0111010101010101;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b0011011100111011;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1101000011111100;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1011111100100000;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b1110100011101000;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b1000100010001000;
    wire [3:0] lut_10_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b0100010111011100;
    wire [3:0] lut_11_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b1111110111011101;
    wire [3:0] lut_12_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b1000111010001000;
    wire [3:0] lut_13_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b1011001010110010;
    wire [3:0] lut_14_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1100110011111110;
    wire [3:0] lut_15_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b1110100011111110;
    wire [3:0] lut_16_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b1110100010000000;
    wire [3:0] lut_17_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b1111111101110001;
    wire [3:0] lut_18_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b0100110101000100;
    wire [3:0] lut_19_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0010000010111111;
    wire [3:0] lut_20_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b1010111100001011;
    wire [3:0] lut_21_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b1011101100100000;
    wire [3:0] lut_22_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0001001001111111;
    wire [3:0] lut_23_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1010001000000000;
    wire [3:0] lut_24_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b1111000101010101;
    wire [3:0] lut_25_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b1100000011110000;
    wire [3:0] lut_26_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1011111100001000;
    wire [3:0] lut_27_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b0000111001001100;
    wire [3:0] lut_28_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b0000000001011111;
    wire [3:0] lut_29_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b0101010111111111;
    wire [3:0] lut_30_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1111110011011100;
    wire [3:0] lut_31_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1111111101000000;
    wire [3:0] lut_32_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b0111000101110001;
    wire [3:0] lut_33_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b0011101100101011;
    wire [3:0] lut_34_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1000000011100000;
    wire [3:0] lut_35_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b0000001100101111;
    wire [3:0] lut_36_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0111000000000000;
    wire [3:0] lut_37_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b1110100011000000;
    wire [3:0] lut_38_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0100000001001100;
    wire [3:0] lut_39_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b0011001100000000;
    wire [3:0] lut_40_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b0010000010101010;
    wire [3:0] lut_41_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b0000111100000000;
    wire [3:0] lut_42_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b1000000010111000;
    wire [3:0] lut_43_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b0000111110111111;
    wire [3:0] lut_44_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b1010101100111111;
    wire [3:0] lut_45_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b0000000011110000;
    wire [3:0] lut_46_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b0000010011001100;
    wire [3:0] lut_47_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b0000011100101111;
    wire [3:0] lut_48_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b0101010111011111;
    wire [3:0] lut_49_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0011000011110000;
    wire [3:0] lut_50_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b0000111000001010;
    wire [3:0] lut_51_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1111011101110000;
    wire [3:0] lut_52_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b1011001010110010;
    wire [3:0] lut_53_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b1011101110111011;
    wire [3:0] lut_54_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b0011101011111111;
    wire [3:0] lut_55_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b0001000100010101;
    wire [3:0] lut_56_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b0000110011101111;
    wire [3:0] lut_57_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b1011101100101011;
    wire [3:0] lut_58_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b0010000010101010;
    wire [3:0] lut_59_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b0101000001110111;
    wire [3:0] lut_60_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b1111001000000000;
    wire [3:0] lut_61_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b1110000011100100;
    wire [3:0] lut_62_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b0101010101010101;
    wire [3:0] lut_63_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b1111111110101010;
    wire [3:0] lut_64_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b1010000011111111;
    wire [3:0] lut_65_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b0000111100011111;
    wire [3:0] lut_66_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b1111110110001101;
    wire [3:0] lut_67_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b0000110001010101;
    wire [3:0] lut_68_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b1101010011110111;
    wire [3:0] lut_69_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b1111001100100010;
    wire [3:0] lut_70_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0101111101011111;
    wire [3:0] lut_71_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b1000111011101111;
    wire [3:0] lut_72_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b0001000001110101;
    wire [3:0] lut_73_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0010000011110010;
    wire [3:0] lut_74_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b1011101100100010;
    wire [3:0] lut_75_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0000000000110011;
    wire [3:0] lut_76_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b1010101000000000;
    wire [3:0] lut_77_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b1111101010111010;
    wire [3:0] lut_78_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b1111111101010101;
    wire [3:0] lut_79_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b1011101011111111;
    wire [3:0] lut_80_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b1110100011111100;
    wire [3:0] lut_81_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1010101110101010;
    wire [3:0] lut_82_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b0011111100111111;
    wire [3:0] lut_83_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b1111101110000010;
    wire [3:0] lut_84_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b1111000010110011;
    wire [3:0] lut_85_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b0100010111110111;
    wire [3:0] lut_86_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b0000000000001101;
    wire [3:0] lut_87_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b0000000000100010;
    wire [3:0] lut_88_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b0001111100010001;
    wire [3:0] lut_89_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1111000010000000;
    wire [3:0] lut_90_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b0000000000001100;
    wire [3:0] lut_91_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1111111101010000;
    wire [3:0] lut_92_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0011011110111111;
    wire [3:0] lut_93_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b0010000010111011;
    wire [3:0] lut_94_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b0010001100111011;
    wire [3:0] lut_95_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1111001100110000;
    wire [3:0] lut_96_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b0000101010101011;
    wire [3:0] lut_97_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1110111011100000;
    wire [3:0] lut_98_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b1111101110111011;
    wire [3:0] lut_99_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1101010011010101;
    wire [3:0] lut_100_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b1111101010101000;
    wire [3:0] lut_101_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b1011001111111111;
    wire [3:0] lut_102_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b0010111110111111;
    wire [3:0] lut_103_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b1010101010000000;
    wire [3:0] lut_104_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1111111110001100;
    wire [3:0] lut_105_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b1100000011110100;
    wire [3:0] lut_106_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b0100110111011101;
    wire [3:0] lut_107_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b0000111111001111;
    wire [3:0] lut_108_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b1110011101100010;
    wire [3:0] lut_109_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b1010000010110111;
    wire [3:0] lut_110_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000000101110111;
    wire [3:0] lut_111_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b1101010011010000;
    wire [3:0] lut_112_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b1111010101010000;
    wire [3:0] lut_113_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1111111111001111;
    wire [3:0] lut_114_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0000000000001100;
    wire [3:0] lut_115_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b1111110101011100;
    wire [3:0] lut_116_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b0000101100001111;
    wire [3:0] lut_117_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1011000011110000;
    wire [3:0] lut_118_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b0010011100000001;
    wire [3:0] lut_119_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b0000101100101011;
    wire [3:0] lut_120_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b1010101010111111;
    wire [3:0] lut_121_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b1100110011101111;
    wire [3:0] lut_122_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b1101110101010101;
    wire [3:0] lut_123_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b0001000101110111;
    wire [3:0] lut_124_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b0001000001110111;
    wire [3:0] lut_125_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b0011011101100111;
    wire [3:0] lut_126_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0111001101110011;
    wire [3:0] lut_127_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b0000110000001101;
    wire [3:0] lut_128_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b0000101000001010;
    wire [3:0] lut_129_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b0011101010101010;
    wire [3:0] lut_130_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b1100000010000000;
    wire [3:0] lut_131_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b1100111000000000;
    wire [3:0] lut_132_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0001000000010010;
    wire [3:0] lut_133_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b0100010001010000;
    wire [3:0] lut_134_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b1111000010111001;
    wire [3:0] lut_135_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b0001010101010111;
    wire [3:0] lut_136_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b1101010101000000;
    wire [3:0] lut_137_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b0111011101010101;
    wire [3:0] lut_138_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b1111110111010100;
    wire [3:0] lut_139_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b0000000001110111;
    wire [3:0] lut_140_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b1110101010000000;
    wire [3:0] lut_141_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b1111101000000000;
    wire [3:0] lut_142_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0000110011101111;
    wire [3:0] lut_143_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b1010100011111110;
    wire [3:0] lut_144_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1110100010000000;
    wire [3:0] lut_145_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1111011101110001;
    wire [3:0] lut_146_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0011000100110000;
    wire [3:0] lut_147_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b1101011101010011;
    wire [3:0] lut_148_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b0101000011010100;
    wire [3:0] lut_149_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b0101010001010101;
    wire [3:0] lut_150_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b0101011101110101;
    wire [3:0] lut_151_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b1110101000000000;
    wire [3:0] lut_152_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1101000101000100;
    wire [3:0] lut_153_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b1100100011011000;
    wire [3:0] lut_154_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b0101111100001100;
    wire [3:0] lut_155_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b0101010111111111;
    wire [3:0] lut_156_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b0010101000101010;
    wire [3:0] lut_157_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b0010000000000111;
    wire [3:0] lut_158_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b0000000000111011;
    wire [3:0] lut_159_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b0000001010100010;
    wire [3:0] lut_160_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b1111100100110000;
    wire [3:0] lut_161_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1011111100101011;
    wire [3:0] lut_162_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b0001111100011111;
    wire [3:0] lut_163_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b1101110011111000;
    wire [3:0] lut_164_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b0010101111111111;
    wire [3:0] lut_165_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b1110101011101010;
    wire [3:0] lut_166_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b0100000001000100;
    wire [3:0] lut_167_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b1000101111111111;
    wire [3:0] lut_168_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b0000000011101110;
    wire [3:0] lut_169_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b1111001011110010;
    wire [3:0] lut_170_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b1000000011001000;
    wire [3:0] lut_171_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b0010101110111111;
    wire [3:0] lut_172_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b1010101100011111;
    wire [3:0] lut_173_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b0000000001110001;
    wire [3:0] lut_174_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1111111111110011;
    wire [3:0] lut_175_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b1010101110111011;
    wire [3:0] lut_176_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b0100010101011111;
    wire [3:0] lut_177_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b0001000011110010;
    wire [3:0] lut_178_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b1011100010111100;
    wire [3:0] lut_179_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b0000100010001110;
    wire [3:0] lut_180_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b1100110100001100;
    wire [3:0] lut_181_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b0000101100000011;
    wire [3:0] lut_182_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b0111000111110111;
    wire [3:0] lut_183_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b0001010100110101;
    wire [3:0] lut_184_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b1010101010101111;
    wire [3:0] lut_185_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b0101010011010100;
    wire [3:0] lut_186_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b1101110110001100;
    wire [3:0] lut_187_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b0100001111000111;
    wire [3:0] lut_188_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b1011001010100000;
    wire [3:0] lut_189_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b1110000011100000;
    wire [3:0] lut_190_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b0111010101010101;
    wire [3:0] lut_191_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b0000110101001111;
    wire [3:0] lut_192_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b0010000011111111;
    wire [3:0] lut_193_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0000111100011111;
    wire [3:0] lut_194_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b1111110111001100;
    wire [3:0] lut_195_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b0001000101110111;
    wire [3:0] lut_196_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b0010101100100010;
    wire [3:0] lut_197_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b1111001010100000;
    wire [3:0] lut_198_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b0101011101000100;
    wire [3:0] lut_199_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b0000111111111111;
    wire [3:0] lut_200_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b1110111010001010;
    wire [3:0] lut_201_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b0010000010110010;
    wire [3:0] lut_202_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b1101010011110001;
    wire [3:0] lut_203_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b0000000000010001;
    wire [3:0] lut_204_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b1101010111111101;
    wire [3:0] lut_205_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b1011101110111010;
    wire [3:0] lut_206_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b0111011100010001;
    wire [3:0] lut_207_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1111010011000000;
    wire [3:0] lut_208_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b0000010100000101;
    wire [3:0] lut_209_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b0000011100001111;
    wire [3:0] lut_210_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b0010111100111111;
    wire [3:0] lut_211_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b1110100011000000;
    wire [3:0] lut_212_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b1100010001000000;
    wire [3:0] lut_213_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1100010111111111;
    wire [3:0] lut_214_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b1111111110110010;
    wire [3:0] lut_215_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b1111111111011100;
    wire [3:0] lut_216_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b1110001011101010;
    wire [3:0] lut_217_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b0000111100111111;
    wire [3:0] lut_218_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b0000000010111011;
    wire [3:0] lut_219_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b0000000000110101;
    wire [3:0] lut_220_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b0101111101001101;
    wire [3:0] lut_221_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b1010100011101100;
    wire [3:0] lut_222_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1110110011101010;
    wire [3:0] lut_223_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b0000100010101010;
    wire [3:0] lut_224_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b1101110101000000;
    wire [3:0] lut_225_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1010001011101011;
    wire [3:0] lut_226_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b0000000001010001;
    wire [3:0] lut_227_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b1111000001110000;
    wire [3:0] lut_228_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b0111000011110011;
    wire [3:0] lut_229_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b0010111111111111;
    wire [3:0] lut_230_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b0011011100111111;
    wire [3:0] lut_231_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b0001111101111111;
    wire [3:0] lut_232_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b0001000101010101;
    wire [3:0] lut_233_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b0100010001110100;
    wire [3:0] lut_234_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b0100110111011101;
    wire [3:0] lut_235_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b1000100011101111;
    wire [3:0] lut_236_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b0111011101110011;
    wire [3:0] lut_237_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b1011111100100011;
    wire [3:0] lut_238_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0000110111011111;
    wire [3:0] lut_239_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b0101010100010011;
    wire [3:0] lut_240_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b0010001000101011;
    wire [3:0] lut_241_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b1111111111001100;
    wire [3:0] lut_242_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b1111111111110011;
    wire [3:0] lut_243_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b1111110101111100;
    wire [3:0] lut_244_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b1100000000000100;
    wire [3:0] lut_245_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b0111001100000000;
    wire [3:0] lut_246_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b0111001100010001;
    wire [3:0] lut_247_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b1110110001001100;
    wire [3:0] lut_248_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b0001011100110011;
    wire [3:0] lut_249_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b1100110111001111;
    wire [3:0] lut_250_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b1101111101011101;
    wire [3:0] lut_251_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b1111111101001110;
    wire [3:0] lut_252_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b1010111010001010;
    wire [3:0] lut_253_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b0111010001010100;
    wire [3:0] lut_254_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b1101110101000101;
    wire [3:0] lut_255_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b1111001101110001;
    wire [3:0] lut_256_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b0000101000001000;
    wire [3:0] lut_257_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b1101000011111000;
    wire [3:0] lut_258_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b0010011000100011;
    wire [3:0] lut_259_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b1100110011010100;
    wire [3:0] lut_260_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b0001000000010000;
    wire [3:0] lut_261_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b0010101110111011;
    wire [3:0] lut_262_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b1111000111111011;
    wire [3:0] lut_263_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b1011111100000000;
    wire [3:0] lut_264_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b1110100011000000;
    wire [3:0] lut_265_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1111111101110111;
    wire [3:0] lut_266_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b0000000011111100;
    wire [3:0] lut_267_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1000101100000010;
    wire [3:0] lut_268_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0000111100001010;
    wire [3:0] lut_269_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b0001100011011101;
    wire [3:0] lut_270_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b1101110000001100;
    wire [3:0] lut_271_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b0101011100000101;
    wire [3:0] lut_272_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b1100000000000000;
    wire [3:0] lut_273_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b1111111101110101;
    wire [3:0] lut_274_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b1110111011001110;
    wire [3:0] lut_275_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b0101011101010111;
    wire [3:0] lut_276_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b1011101100000010;
    wire [3:0] lut_277_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b0101010001010000;
    wire [3:0] lut_278_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b1110101100000011;
    wire [3:0] lut_279_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b0001111100111111;
    wire [3:0] lut_280_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b0010001100110111;
    wire [3:0] lut_281_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b1011101010100000;
    wire [3:0] lut_282_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b0000001111110111;
    wire [3:0] lut_283_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b1100101010000000;
    wire [3:0] lut_284_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b0000101000001010;
    wire [3:0] lut_285_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b0010000100000111;
    wire [3:0] lut_286_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b0010001000101010;
    wire [3:0] lut_287_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b1101110111011101;
    wire [3:0] lut_288_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b0000011101011111;
    wire [3:0] lut_289_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b1011101100101011;
    wire [3:0] lut_290_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b0111111100011111;
    wire [3:0] lut_291_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b0001000101110001;
    wire [3:0] lut_292_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b0000111111111111;
    wire [3:0] lut_293_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1110100011000000;
    wire [3:0] lut_294_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b1111110011110100;
    wire [3:0] lut_295_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b1000101111111111;
    wire [3:0] lut_296_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b0111111100010001;
    wire [3:0] lut_297_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b0000110101001100;
    wire [3:0] lut_298_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b1000000011101000;
    wire [3:0] lut_299_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b1111010101010000;
    wire [3:0] lut_300_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b0101010011100000;
    wire [3:0] lut_301_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b1011000001110000;
    wire [3:0] lut_302_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b1100110111001101;
    wire [3:0] lut_303_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b1101010011000100;
    wire [3:0] lut_304_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b1011001000100000;
    wire [3:0] lut_305_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b0011000101110011;
    wire [3:0] lut_306_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b0100001111110011;
    wire [3:0] lut_307_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b0101110001011110;
    wire [3:0] lut_308_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b1100111100001100;
    wire [3:0] lut_309_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b1011111100111011;
    wire [3:0] lut_310_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b1111000111110011;
    wire [3:0] lut_311_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1111111111101110;
    wire [3:0] lut_312_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b0010111010101111;
    wire [3:0] lut_313_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b0010111100001011;
    wire [3:0] lut_314_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b0000111100000100;
    wire [3:0] lut_315_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b0001000111110111;
    wire [3:0] lut_316_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b1011101010100000;
    wire [3:0] lut_317_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0001101101010101;
    wire [3:0] lut_318_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b1100111010001110;
    wire [3:0] lut_319_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b1110111010101111;
    wire [3:0] lut_320_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0010001111111011;
    wire [3:0] lut_321_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b0101011100010011;
    wire [3:0] lut_322_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b1111111111001100;
    wire [3:0] lut_323_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b1110111110001110;
    wire [3:0] lut_324_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b1101000011110000;
    wire [3:0] lut_325_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b1110110011111100;
    wire [3:0] lut_326_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b1110000010100100;
    wire [3:0] lut_327_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b1000101010101111;
    wire [3:0] lut_328_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b1111001111110011;
    wire [3:0] lut_329_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b1111111111000000;
    wire [3:0] lut_330_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b0100010011111101;
    wire [3:0] lut_331_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b0000000000010001;
    wire [3:0] lut_332_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b0101010111111111;
    wire [3:0] lut_333_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b0000010011000101;
    wire [3:0] lut_334_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0011111100101111;
    wire [3:0] lut_335_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b0000101100001001;
    wire [3:0] lut_336_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b0000010011101111;
    wire [3:0] lut_337_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b0000010001111111;
    wire [3:0] lut_338_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b1101000011110000;
    wire [3:0] lut_339_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b1111110111000000;
    wire [3:0] lut_340_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b1101110001000000;
    wire [3:0] lut_341_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b0001000001110011;
    wire [3:0] lut_342_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b1101010111110000;
    wire [3:0] lut_343_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1111110111111100;
    wire [3:0] lut_344_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b0001111100010001;
    wire [3:0] lut_345_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b1111100000000000;
    wire [3:0] lut_346_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b0000000000111010;
    wire [3:0] lut_347_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0000000000100101;
    wire [3:0] lut_348_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b1100110000000100;
    wire [3:0] lut_349_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b1010111111111101;
    wire [3:0] lut_350_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b1111101110110000;
    wire [3:0] lut_351_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b1111010101110101;
    wire [3:0] lut_352_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b1111000001110011;
    wire [3:0] lut_353_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b1000100010001100;
    wire [3:0] lut_354_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b1111001111110011;
    wire [3:0] lut_355_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b1100010011001100;
    wire [3:0] lut_356_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b0000010101010111;
    wire [3:0] lut_357_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b0101110000000000;
    wire [3:0] lut_358_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b0010111110111111;
    wire [3:0] lut_359_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b1000101010001110;
    wire [3:0] lut_360_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b1110111100000000;
    wire [3:0] lut_361_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b1101010011011100;
    wire [3:0] lut_362_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b1111001100110000;
    wire [3:0] lut_363_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b0000100011101111;
    wire [3:0] lut_364_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b1000110011001111;
    wire [3:0] lut_365_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b0000110010001101;
    wire [3:0] lut_366_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b0001111101111111;
    wire [3:0] lut_367_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b1100111110001000;
    wire [3:0] lut_368_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b1101110111011100;
    wire [3:0] lut_369_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b0010001010111011;
    wire [3:0] lut_370_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b0000000000001100;
    wire [3:0] lut_371_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b1111110011111110;
    wire [3:0] lut_372_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b0010111000100111;
    wire [3:0] lut_373_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b1110110011111101;
    wire [3:0] lut_374_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b0111000100010001;
    wire [3:0] lut_375_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b1010101110001011;
    wire [3:0] lut_376_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b1101010111000000;
    wire [3:0] lut_377_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b1100111011101110;
    wire [3:0] lut_378_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1111000011110111;
    wire [3:0] lut_379_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b1110000010110011;
    wire [3:0] lut_380_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b0101000001110111;
    wire [3:0] lut_381_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b0000100010001100;
    wire [3:0] lut_382_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b0011000010110011;
    wire [3:0] lut_383_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0000110000001111;
    wire [3:0] lut_384_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b1000111000001010;
    wire [3:0] lut_385_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b1011100110111111;
    wire [3:0] lut_386_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b1101000010001000;
    wire [3:0] lut_387_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b0101010111110101;
    wire [3:0] lut_388_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b1111010101000100;
    wire [3:0] lut_389_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b1110001001000000;
    wire [3:0] lut_390_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b0000011100000100;
    wire [3:0] lut_391_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b1011101110100000;
    wire [3:0] lut_392_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b1101010000000000;
    wire [3:0] lut_393_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b0111111101110111;
    wire [3:0] lut_394_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b1111111101010001;
    wire [3:0] lut_395_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b0000001100001011;
    wire [3:0] lut_396_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b1010111000001000;
    wire [3:0] lut_397_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b0010101010111010;
    wire [3:0] lut_398_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b0111001101010001;
    wire [3:0] lut_399_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b1010101010111011;
    wire [3:0] lut_400_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b1110100010000000;
    wire [3:0] lut_401_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b0000100010001010;
    wire [3:0] lut_402_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b0001000000110000;
    wire [3:0] lut_403_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b0010000010111111;
    wire [3:0] lut_404_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b1010111100001011;
    wire [3:0] lut_405_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0100010001010111;
    wire [3:0] lut_406_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b0000001100000001;
    wire [3:0] lut_407_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b1110010001010101;
    wire [3:0] lut_408_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b0000101100111111;
    wire [3:0] lut_409_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b1011111100001011;
    wire [3:0] lut_410_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b0100000111001011;
    wire [3:0] lut_411_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b0011000011111011;
    wire [3:0] lut_412_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b0011001100001011;
    wire [3:0] lut_413_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0010000100000111;
    wire [3:0] lut_414_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b0000100100001011;
    wire [3:0] lut_415_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b0011000010111011;
    wire [3:0] lut_416_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b0000110010001110;
    wire [3:0] lut_417_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b1010101100111011;
    wire [3:0] lut_418_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b0111111100011111;
    wire [3:0] lut_419_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b1000100010001010;
    wire [3:0] lut_420_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b0010101111111111;
    wire [3:0] lut_421_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b1010101010101000;
    wire [3:0] lut_422_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b1111110011111100;
    wire [3:0] lut_423_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b0000111111011111;
    wire [3:0] lut_424_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b0000000011101110;
    wire [3:0] lut_425_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b0100110100001101;
    wire [3:0] lut_426_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b1000000010101000;
    wire [3:0] lut_427_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b1101010101000100;
    wire [3:0] lut_428_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b0111000011100000;
    wire [3:0] lut_429_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b1011000010110000;
    wire [3:0] lut_430_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b1111011101010000;
    wire [3:0] lut_431_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b1000101011101011;
    wire [3:0] lut_432_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b1011001010100010;
    wire [3:0] lut_433_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b1110111100101111;
    wire [3:0] lut_434_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b1000111000001011;
    wire [3:0] lut_435_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b1111111101110000;
    wire [3:0] lut_436_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b0100110100000000;
    wire [3:0] lut_437_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b0000000001000100;
    wire [3:0] lut_438_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b1111010110110011;
    wire [3:0] lut_439_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b1110110011001110;
    wire [3:0] lut_440_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b1000110011001110;
    wire [3:0] lut_441_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b0011101100101011;
    wire [3:0] lut_442_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1110110110001101;
    wire [3:0] lut_443_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b1111010011000000;
    wire [3:0] lut_444_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b1011101000100010;
    wire [3:0] lut_445_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b1111000011111010;
    wire [3:0] lut_446_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b0100111011001110;
    wire [3:0] lut_447_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b0001111100101111;
    wire [3:0] lut_448_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b0010001110110011;
    wire [3:0] lut_449_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b0011011100110011;
    wire [3:0] lut_450_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b1110000010000010;
    wire [3:0] lut_451_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b1111111110101110;
    wire [3:0] lut_452_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b0010001000100010;
    wire [3:0] lut_453_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0001111100011101;
    wire [3:0] lut_454_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b0010000001100100;
    wire [3:0] lut_455_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b0010111111111111;
    wire [3:0] lut_456_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b1111111110110010;
    wire [3:0] lut_457_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b0110000001110010;
    wire [3:0] lut_458_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b0101010011111101;
    wire [3:0] lut_459_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b0000000100000101;
    wire [3:0] lut_460_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b1110111000001000;
    wire [3:0] lut_461_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b1101101000001010;
    wire [3:0] lut_462_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b1111010100000000;
    wire [3:0] lut_463_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b1110101011101110;
    wire [3:0] lut_464_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b0001010100000001;
    wire [3:0] lut_465_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b1010101100000000;
    wire [3:0] lut_466_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1011101110100010;
    wire [3:0] lut_467_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b1101111111010100;
    wire [3:0] lut_468_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b1010101010101011;
    wire [3:0] lut_469_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b0100010111111111;
    wire [3:0] lut_470_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b0000101000001111;
    wire [3:0] lut_471_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b0000001000100011;
    wire [3:0] lut_472_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b1111000011111111;
    wire [3:0] lut_473_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b1111111010000000;
    wire [3:0] lut_474_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b0000000000111110;
    wire [3:0] lut_475_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b1111110111011000;
    wire [3:0] lut_476_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b0101111101011101;
    wire [3:0] lut_477_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b0111010100010000;
    wire [3:0] lut_478_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b1111111011000000;
    wire [3:0] lut_479_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b1111011101110101;
    wire [3:0] lut_480_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b1111100011010000;
    wire [3:0] lut_481_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b1101111100000101;
    wire [3:0] lut_482_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b0000110000001100;
    wire [3:0] lut_483_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b1101000011010100;
    wire [3:0] lut_484_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b0111000011110011;
    wire [3:0] lut_485_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b1011000011110000;
    wire [3:0] lut_486_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b0010111110111111;
    wire [3:0] lut_487_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1100111010001010;
    wire [3:0] lut_488_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b1110111011001010;
    wire [3:0] lut_489_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b1010111100001111;
    wire [3:0] lut_490_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b0011001100110011;
    wire [3:0] lut_491_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b1111000000010000;
    wire [3:0] lut_492_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b0111011101110011;
    wire [3:0] lut_493_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b1000110010101111;
    wire [3:0] lut_494_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b1110110000000000;
    wire [3:0] lut_495_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b1110000011110000;
    wire [3:0] lut_496_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b0000001011101010;
    wire [3:0] lut_497_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b0000100000111001;
    wire [3:0] lut_498_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b0000010000001100;
    wire [3:0] lut_499_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b1111110001011100;
    wire [3:0] lut_500_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b1110111100001000;
    wire [3:0] lut_501_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b0001011100000010;
    wire [3:0] lut_502_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b1000101010001110;
    wire [3:0] lut_503_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b1111110100100100;
    wire [3:0] lut_504_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b0000000011101010;
    wire [3:0] lut_505_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b1111000100010000;
    wire [3:0] lut_506_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b0001111100001101;
    wire [3:0] lut_507_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b1110111000001000;
    wire [3:0] lut_508_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b1100111100000000;
    wire [3:0] lut_509_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b1000110011001000;
    wire [3:0] lut_510_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0011000011111011;
    wire [3:0] lut_511_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [15:0] lut_512_table = 16'b0000110011001110;
    wire [3:0] lut_512_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [15:0] lut_513_table = 16'b0111000111110111;
    wire [3:0] lut_513_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [15:0] lut_514_table = 16'b0010111111100110;
    wire [3:0] lut_514_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [15:0] lut_515_table = 16'b1100110001001101;
    wire [3:0] lut_515_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [15:0] lut_516_table = 16'b0010101000001010;
    wire [3:0] lut_516_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [15:0] lut_517_table = 16'b1010111011101111;
    wire [3:0] lut_517_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [15:0] lut_518_table = 16'b1100001001000000;
    wire [3:0] lut_518_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [15:0] lut_519_table = 16'b1111000010111000;
    wire [3:0] lut_519_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [15:0] lut_520_table = 16'b0011101100100011;
    wire [3:0] lut_520_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [15:0] lut_521_table = 16'b1111100011100000;
    wire [3:0] lut_521_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [15:0] lut_522_table = 16'b1000000011001000;
    wire [3:0] lut_522_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [15:0] lut_523_table = 16'b0010001000101010;
    wire [3:0] lut_523_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [15:0] lut_524_table = 16'b1101010011110101;
    wire [3:0] lut_524_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [15:0] lut_525_table = 16'b0101010101110111;
    wire [3:0] lut_525_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [15:0] lut_526_table = 16'b0101010101010101;
    wire [3:0] lut_526_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [15:0] lut_527_table = 16'b1110011001110011;
    wire [3:0] lut_527_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [15:0] lut_528_table = 16'b0001001100010000;
    wire [3:0] lut_528_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [15:0] lut_529_table = 16'b1111101010100000;
    wire [3:0] lut_529_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [15:0] lut_530_table = 16'b0000100010001110;
    wire [3:0] lut_530_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [15:0] lut_531_table = 16'b1110111110101111;
    wire [3:0] lut_531_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [15:0] lut_532_table = 16'b1101011101000001;
    wire [3:0] lut_532_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [15:0] lut_533_table = 16'b0101010101010101;
    wire [3:0] lut_533_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [15:0] lut_534_table = 16'b1010101100101011;
    wire [3:0] lut_534_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [15:0] lut_535_table = 16'b1110000011101010;
    wire [3:0] lut_535_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [15:0] lut_536_table = 16'b1011001000000000;
    wire [3:0] lut_536_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [15:0] lut_537_table = 16'b0000111110111011;
    wire [3:0] lut_537_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [15:0] lut_538_table = 16'b0011011100000111;
    wire [3:0] lut_538_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [15:0] lut_539_table = 16'b0011111000101000;
    wire [3:0] lut_539_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [15:0] lut_540_table = 16'b0001111101111111;
    wire [3:0] lut_540_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [15:0] lut_541_table = 16'b0000101000001010;
    wire [3:0] lut_541_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [15:0] lut_542_table = 16'b0101110111111111;
    wire [3:0] lut_542_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [15:0] lut_543_table = 16'b1111111111011100;
    wire [3:0] lut_543_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [15:0] lut_544_table = 16'b1111110101011101;
    wire [3:0] lut_544_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [15:0] lut_545_table = 16'b0000010011101111;
    wire [3:0] lut_545_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [15:0] lut_546_table = 16'b0100000011010100;
    wire [3:0] lut_546_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [15:0] lut_547_table = 16'b0101111100001111;
    wire [3:0] lut_547_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [15:0] lut_548_table = 16'b0011000101110001;
    wire [3:0] lut_548_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [15:0] lut_549_table = 16'b0010101111111111;
    wire [3:0] lut_549_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [15:0] lut_550_table = 16'b0001111100001111;
    wire [3:0] lut_550_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [15:0] lut_551_table = 16'b1111111010101000;
    wire [3:0] lut_551_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [15:0] lut_552_table = 16'b1100111011111111;
    wire [3:0] lut_552_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [15:0] lut_553_table = 16'b0011001110111010;
    wire [3:0] lut_553_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [15:0] lut_554_table = 16'b0100110101001100;
    wire [3:0] lut_554_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [15:0] lut_555_table = 16'b1000000011100000;
    wire [3:0] lut_555_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [15:0] lut_556_table = 16'b1111110111010100;
    wire [3:0] lut_556_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [15:0] lut_557_table = 16'b1010111100101010;
    wire [3:0] lut_557_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [15:0] lut_558_table = 16'b0000000001110001;
    wire [3:0] lut_558_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [15:0] lut_559_table = 16'b1100110111001101;
    wire [3:0] lut_559_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [15:0] lut_560_table = 16'b1111110000000000;
    wire [3:0] lut_560_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [15:0] lut_561_table = 16'b1010001010100000;
    wire [3:0] lut_561_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [15:0] lut_562_table = 16'b0100111100001111;
    wire [3:0] lut_562_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [15:0] lut_563_table = 16'b1111100011111100;
    wire [3:0] lut_563_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [15:0] lut_564_table = 16'b1111010101110000;
    wire [3:0] lut_564_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [15:0] lut_565_table = 16'b1011001011110010;
    wire [3:0] lut_565_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [15:0] lut_566_table = 16'b0000000001010101;
    wire [3:0] lut_566_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [15:0] lut_567_table = 16'b1111000100110011;
    wire [3:0] lut_567_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [15:0] lut_568_table = 16'b1110111011001110;
    wire [3:0] lut_568_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [15:0] lut_569_table = 16'b0010001011101111;
    wire [3:0] lut_569_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [15:0] lut_570_table = 16'b0100000011111111;
    wire [3:0] lut_570_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [15:0] lut_571_table = 16'b0001011100000101;
    wire [3:0] lut_571_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [15:0] lut_572_table = 16'b0000101000111111;
    wire [3:0] lut_572_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [15:0] lut_573_table = 16'b1011101010100000;
    wire [3:0] lut_573_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [15:0] lut_574_table = 16'b0000111001010101;
    wire [3:0] lut_574_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [15:0] lut_575_table = 16'b1111010101010000;
    wire [3:0] lut_575_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [15:0] lut_576_table = 16'b0100000001010100;
    wire [3:0] lut_576_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [15:0] lut_577_table = 16'b0010001011111011;
    wire [3:0] lut_577_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [15:0] lut_578_table = 16'b0000101000001111;
    wire [3:0] lut_578_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [15:0] lut_579_table = 16'b0101111101001101;
    wire [3:0] lut_579_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [15:0] lut_580_table = 16'b0001000001110001;
    wire [3:0] lut_580_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [15:0] lut_581_table = 16'b1101110011011101;
    wire [3:0] lut_581_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [15:0] lut_582_table = 16'b0000111100010111;
    wire [3:0] lut_582_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [15:0] lut_583_table = 16'b0010000001110100;
    wire [3:0] lut_583_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [15:0] lut_584_table = 16'b0111000101010000;
    wire [3:0] lut_584_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [15:0] lut_585_table = 16'b1111011111110011;
    wire [3:0] lut_585_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [15:0] lut_586_table = 16'b1101111111001101;
    wire [3:0] lut_586_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [15:0] lut_587_table = 16'b0010101100000010;
    wire [3:0] lut_587_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [15:0] lut_588_table = 16'b0000110100000001;
    wire [3:0] lut_588_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [15:0] lut_589_table = 16'b0101010111110101;
    wire [3:0] lut_589_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [15:0] lut_590_table = 16'b1101101100001000;
    wire [3:0] lut_590_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [15:0] lut_591_table = 16'b0001010110001100;
    wire [3:0] lut_591_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [15:0] lut_592_table = 16'b1000000011000100;
    wire [3:0] lut_592_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [15:0] lut_593_table = 16'b1111111100000000;
    wire [3:0] lut_593_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [15:0] lut_594_table = 16'b0101010001110111;
    wire [3:0] lut_594_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [15:0] lut_595_table = 16'b0101000011111101;
    wire [3:0] lut_595_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [15:0] lut_596_table = 16'b0000001100111111;
    wire [3:0] lut_596_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [15:0] lut_597_table = 16'b0011101111111111;
    wire [3:0] lut_597_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [15:0] lut_598_table = 16'b0001000001110001;
    wire [3:0] lut_598_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [15:0] lut_599_table = 16'b0000000001001111;
    wire [3:0] lut_599_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [15:0] lut_600_table = 16'b1101110111110100;
    wire [3:0] lut_600_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [15:0] lut_601_table = 16'b0000111100011000;
    wire [3:0] lut_601_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [15:0] lut_602_table = 16'b0101010001010100;
    wire [3:0] lut_602_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [15:0] lut_603_table = 16'b0000100010111011;
    wire [3:0] lut_603_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [15:0] lut_604_table = 16'b0010001000100111;
    wire [3:0] lut_604_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [15:0] lut_605_table = 16'b1010000010100000;
    wire [3:0] lut_605_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [15:0] lut_606_table = 16'b1011110111101100;
    wire [3:0] lut_606_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [15:0] lut_607_table = 16'b1111111011110000;
    wire [3:0] lut_607_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [15:0] lut_608_table = 16'b1000101010001010;
    wire [3:0] lut_608_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [15:0] lut_609_table = 16'b1000111010101011;
    wire [3:0] lut_609_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [15:0] lut_610_table = 16'b0010001010101110;
    wire [3:0] lut_610_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [15:0] lut_611_table = 16'b1100111110001110;
    wire [3:0] lut_611_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [15:0] lut_612_table = 16'b0011001100110011;
    wire [3:0] lut_612_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [15:0] lut_613_table = 16'b0001000001110101;
    wire [3:0] lut_613_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [15:0] lut_614_table = 16'b1010101011111011;
    wire [3:0] lut_614_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [15:0] lut_615_table = 16'b1101010100000000;
    wire [3:0] lut_615_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [15:0] lut_616_table = 16'b0111011101110111;
    wire [3:0] lut_616_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [15:0] lut_617_table = 16'b0101111100000100;
    wire [3:0] lut_617_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [15:0] lut_618_table = 16'b0100010011110100;
    wire [3:0] lut_618_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [15:0] lut_619_table = 16'b1011001000000000;
    wire [3:0] lut_619_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [15:0] lut_620_table = 16'b1000110011101111;
    wire [3:0] lut_620_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [15:0] lut_621_table = 16'b0111001100110000;
    wire [3:0] lut_621_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [15:0] lut_622_table = 16'b0000001100000101;
    wire [3:0] lut_622_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [15:0] lut_623_table = 16'b0001011101011111;
    wire [3:0] lut_623_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [15:0] lut_624_table = 16'b0000100000101110;
    wire [3:0] lut_624_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [15:0] lut_625_table = 16'b1010101010101010;
    wire [3:0] lut_625_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [15:0] lut_626_table = 16'b1111010101010101;
    wire [3:0] lut_626_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [15:0] lut_627_table = 16'b0000000000001100;
    wire [3:0] lut_627_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [15:0] lut_628_table = 16'b0000001000100011;
    wire [3:0] lut_628_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [15:0] lut_629_table = 16'b1110011000000101;
    wire [3:0] lut_629_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [15:0] lut_630_table = 16'b1100110011111111;
    wire [3:0] lut_630_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [15:0] lut_631_table = 16'b1010111110001000;
    wire [3:0] lut_631_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [15:0] lut_632_table = 16'b0000001001110011;
    wire [3:0] lut_632_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [15:0] lut_633_table = 16'b0010101000111111;
    wire [3:0] lut_633_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [15:0] lut_634_table = 16'b0000111011101111;
    wire [3:0] lut_634_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [15:0] lut_635_table = 16'b0100111100001101;
    wire [3:0] lut_635_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [15:0] lut_636_table = 16'b1110101010001000;
    wire [3:0] lut_636_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [15:0] lut_637_table = 16'b1100111110001000;
    wire [3:0] lut_637_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [15:0] lut_638_table = 16'b1110011100010111;
    wire [3:0] lut_638_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [15:0] lut_639_table = 16'b0000101010101010;
    wire [3:0] lut_639_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub3
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        639:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        639:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub3_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub3_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub3_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [639:0]  in_data,
            output wire [639:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1100110011101111;
    wire [3:0] lut_0_select = {
                             in_data[459],
                             in_data[432],
                             in_data[227],
                             in_data[285]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b1101010111010101;
    wire [3:0] lut_1_select = {
                             in_data[4],
                             in_data[246],
                             in_data[502],
                             in_data[312]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b0011001100010000;
    wire [3:0] lut_2_select = {
                             in_data[638],
                             in_data[287],
                             in_data[633],
                             in_data[148]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1101010100000000;
    wire [3:0] lut_3_select = {
                             in_data[507],
                             in_data[175],
                             in_data[521],
                             in_data[590]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b1100111100001100;
    wire [3:0] lut_4_select = {
                             in_data[413],
                             in_data[153],
                             in_data[196],
                             in_data[123]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b0000111100001010;
    wire [3:0] lut_5_select = {
                             in_data[99],
                             in_data[212],
                             in_data[608],
                             in_data[105]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b1010101000000000;
    wire [3:0] lut_6_select = {
                             in_data[71],
                             in_data[252],
                             in_data[98],
                             in_data[551]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1101110001000000;
    wire [3:0] lut_7_select = {
                             in_data[357],
                             in_data[43],
                             in_data[419],
                             in_data[199]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1111110110000000;
    wire [3:0] lut_8_select = {
                             in_data[606],
                             in_data[247],
                             in_data[472],
                             in_data[19]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b0101000101110001;
    wire [3:0] lut_9_select = {
                             in_data[211],
                             in_data[586],
                             in_data[163],
                             in_data[433]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b0010111100110111;
    wire [3:0] lut_10_select = {
                             in_data[569],
                             in_data[381],
                             in_data[441],
                             in_data[429]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b1111001011110010;
    wire [3:0] lut_11_select = {
                             in_data[282],
                             in_data[438],
                             in_data[360],
                             in_data[113]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b1000000011111110;
    wire [3:0] lut_12_select = {
                             in_data[207],
                             in_data[451],
                             in_data[359],
                             in_data[585]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0100010100010101;
    wire [3:0] lut_13_select = {
                             in_data[155],
                             in_data[293],
                             in_data[573],
                             in_data[42]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0011001101110000;
    wire [3:0] lut_14_select = {
                             in_data[25],
                             in_data[146],
                             in_data[292],
                             in_data[192]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1000111010101010;
    wire [3:0] lut_15_select = {
                             in_data[92],
                             in_data[388],
                             in_data[603],
                             in_data[430]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b0011101100110011;
    wire [3:0] lut_16_select = {
                             in_data[93],
                             in_data[575],
                             in_data[464],
                             in_data[232]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b1111110101010100;
    wire [3:0] lut_17_select = {
                             in_data[520],
                             in_data[300],
                             in_data[107],
                             in_data[504]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b1101010011111101;
    wire [3:0] lut_18_select = {
                             in_data[242],
                             in_data[161],
                             in_data[533],
                             in_data[324]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b0100000011110000;
    wire [3:0] lut_19_select = {
                             in_data[129],
                             in_data[594],
                             in_data[330],
                             in_data[114]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0111111100010001;
    wire [3:0] lut_20_select = {
                             in_data[144],
                             in_data[637],
                             in_data[343],
                             in_data[183]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b1100000111000001;
    wire [3:0] lut_21_select = {
                             in_data[185],
                             in_data[191],
                             in_data[170],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b1110110011111111;
    wire [3:0] lut_22_select = {
                             in_data[344],
                             in_data[220],
                             in_data[371],
                             in_data[261]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0001000101011111;
    wire [3:0] lut_23_select = {
                             in_data[409],
                             in_data[178],
                             in_data[281],
                             in_data[498]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b0111000001000000;
    wire [3:0] lut_24_select = {
                             in_data[34],
                             in_data[122],
                             in_data[214],
                             in_data[505]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0011001100110011;
    wire [3:0] lut_25_select = {
                             in_data[296],
                             in_data[591],
                             in_data[598],
                             in_data[424]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b0111000001110100;
    wire [3:0] lut_26_select = {
                             in_data[313],
                             in_data[154],
                             in_data[530],
                             in_data[570]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1110101110101010;
    wire [3:0] lut_27_select = {
                             in_data[222],
                             in_data[609],
                             in_data[280],
                             in_data[66]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b0101111100001100;
    wire [3:0] lut_28_select = {
                             in_data[83],
                             in_data[494],
                             in_data[140],
                             in_data[69]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b0011001100110011;
    wire [3:0] lut_29_select = {
                             in_data[37],
                             in_data[180],
                             in_data[600],
                             in_data[532]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b0100010101001101;
    wire [3:0] lut_30_select = {
                             in_data[40],
                             in_data[514],
                             in_data[64],
                             in_data[453]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1110000011111111;
    wire [3:0] lut_31_select = {
                             in_data[310],
                             in_data[230],
                             in_data[528],
                             in_data[455]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1110111100001111;
    wire [3:0] lut_32_select = {
                             in_data[583],
                             in_data[260],
                             in_data[560],
                             in_data[412]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b1101111011001100;
    wire [3:0] lut_33_select = {
                             in_data[24],
                             in_data[461],
                             in_data[68],
                             in_data[82]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1010101010101010;
    wire [3:0] lut_34_select = {
                             in_data[350],
                             in_data[307],
                             in_data[120],
                             in_data[20]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1100110011001100;
    wire [3:0] lut_35_select = {
                             in_data[554],
                             in_data[632],
                             in_data[595],
                             in_data[563]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b1101111101011101;
    wire [3:0] lut_36_select = {
                             in_data[431],
                             in_data[386],
                             in_data[354],
                             in_data[164]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0011111011111010;
    wire [3:0] lut_37_select = {
                             in_data[284],
                             in_data[512],
                             in_data[139],
                             in_data[26]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b1011111100001010;
    wire [3:0] lut_38_select = {
                             in_data[204],
                             in_data[380],
                             in_data[465],
                             in_data[210]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0000101100010111;
    wire [3:0] lut_39_select = {
                             in_data[397],
                             in_data[390],
                             in_data[97],
                             in_data[221]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b0011101100001111;
    wire [3:0] lut_40_select = {
                             in_data[198],
                             in_data[500],
                             in_data[104],
                             in_data[422]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b1111000001110001;
    wire [3:0] lut_41_select = {
                             in_data[151],
                             in_data[63],
                             in_data[538],
                             in_data[111]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b1111111100001000;
    wire [3:0] lut_42_select = {
                             in_data[336],
                             in_data[171],
                             in_data[395],
                             in_data[270]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0010001000001010;
    wire [3:0] lut_43_select = {
                             in_data[11],
                             in_data[169],
                             in_data[301],
                             in_data[394]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b1111111110001100;
    wire [3:0] lut_44_select = {
                             in_data[50],
                             in_data[478],
                             in_data[233],
                             in_data[264]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b1111010011010000;
    wire [3:0] lut_45_select = {
                             in_data[238],
                             in_data[321],
                             in_data[138],
                             in_data[486]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b1111010000000000;
    wire [3:0] lut_46_select = {
                             in_data[450],
                             in_data[434],
                             in_data[517],
                             in_data[546]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b1110000010100000;
    wire [3:0] lut_47_select = {
                             in_data[9],
                             in_data[1],
                             in_data[383],
                             in_data[278]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b1100100011101111;
    wire [3:0] lut_48_select = {
                             in_data[224],
                             in_data[249],
                             in_data[414],
                             in_data[579]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b1110000001000000;
    wire [3:0] lut_49_select = {
                             in_data[187],
                             in_data[543],
                             in_data[124],
                             in_data[541]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0000000001010111;
    wire [3:0] lut_50_select = {
                             in_data[518],
                             in_data[197],
                             in_data[471],
                             in_data[561]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b1111101010101000;
    wire [3:0] lut_51_select = {
                             in_data[240],
                             in_data[589],
                             in_data[635],
                             in_data[341]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1000100010110000;
    wire [3:0] lut_52_select = {
                             in_data[411],
                             in_data[30],
                             in_data[447],
                             in_data[339]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b1100010001010101;
    wire [3:0] lut_53_select = {
                             in_data[477],
                             in_data[147],
                             in_data[338],
                             in_data[62]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b1111111111111010;
    wire [3:0] lut_54_select = {
                             in_data[580],
                             in_data[346],
                             in_data[168],
                             in_data[203]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b1111111100101010;
    wire [3:0] lut_55_select = {
                             in_data[558],
                             in_data[226],
                             in_data[487],
                             in_data[488]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b1111001100110010;
    wire [3:0] lut_56_select = {
                             in_data[5],
                             in_data[298],
                             in_data[127],
                             in_data[476]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b1111101011111010;
    wire [3:0] lut_57_select = {
                             in_data[454],
                             in_data[315],
                             in_data[448],
                             in_data[27]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b1111010111110000;
    wire [3:0] lut_58_select = {
                             in_data[463],
                             in_data[65],
                             in_data[536],
                             in_data[255]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b1010111110101111;
    wire [3:0] lut_59_select = {
                             in_data[160],
                             in_data[45],
                             in_data[392],
                             in_data[539]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b1111010101110000;
    wire [3:0] lut_60_select = {
                             in_data[28],
                             in_data[391],
                             in_data[529],
                             in_data[218]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b1011111100100011;
    wire [3:0] lut_61_select = {
                             in_data[345],
                             in_data[581],
                             in_data[557],
                             in_data[481]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b1100000011111000;
    wire [3:0] lut_62_select = {
                             in_data[480],
                             in_data[425],
                             in_data[250],
                             in_data[396]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b1010001011111011;
    wire [3:0] lut_63_select = {
                             in_data[248],
                             in_data[58],
                             in_data[545],
                             in_data[624]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b0000110010001101;
    wire [3:0] lut_64_select = {
                             in_data[70],
                             in_data[88],
                             in_data[442],
                             in_data[439]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b1000111010001010;
    wire [3:0] lut_65_select = {
                             in_data[437],
                             in_data[95],
                             in_data[17],
                             in_data[382]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b1110000011100000;
    wire [3:0] lut_66_select = {
                             in_data[564],
                             in_data[179],
                             in_data[121],
                             in_data[510]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b0000111100000011;
    wire [3:0] lut_67_select = {
                             in_data[7],
                             in_data[59],
                             in_data[332],
                             in_data[374]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b0111000101110011;
    wire [3:0] lut_68_select = {
                             in_data[491],
                             in_data[402],
                             in_data[616],
                             in_data[614]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b1111111100100010;
    wire [3:0] lut_69_select = {
                             in_data[254],
                             in_data[209],
                             in_data[446],
                             in_data[239]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b0101010001000100;
    wire [3:0] lut_70_select = {
                             in_data[599],
                             in_data[256],
                             in_data[231],
                             in_data[547]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0101011101011111;
    wire [3:0] lut_71_select = {
                             in_data[612],
                             in_data[152],
                             in_data[410],
                             in_data[368]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b1111111100001101;
    wire [3:0] lut_72_select = {
                             in_data[131],
                             in_data[143],
                             in_data[316],
                             in_data[35]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b1011101100100010;
    wire [3:0] lut_73_select = {
                             in_data[277],
                             in_data[13],
                             in_data[337],
                             in_data[184]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b1010000010110000;
    wire [3:0] lut_74_select = {
                             in_data[400],
                             in_data[12],
                             in_data[605],
                             in_data[349]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b0010001000100010;
    wire [3:0] lut_75_select = {
                             in_data[23],
                             in_data[362],
                             in_data[162],
                             in_data[537]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0101110001000000;
    wire [3:0] lut_76_select = {
                             in_data[376],
                             in_data[94],
                             in_data[331],
                             in_data[492]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b1101010100000000;
    wire [3:0] lut_77_select = {
                             in_data[286],
                             in_data[55],
                             in_data[358],
                             in_data[257]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b1111101011110011;
    wire [3:0] lut_78_select = {
                             in_data[513],
                             in_data[39],
                             in_data[617],
                             in_data[565]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b1010111100001111;
    wire [3:0] lut_79_select = {
                             in_data[577],
                             in_data[290],
                             in_data[452],
                             in_data[630]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b1111010011110101;
    wire [3:0] lut_80_select = {
                             in_data[615],
                             in_data[87],
                             in_data[351],
                             in_data[302]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b0101011101110111;
    wire [3:0] lut_81_select = {
                             in_data[370],
                             in_data[550],
                             in_data[172],
                             in_data[493]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1101010111010101;
    wire [3:0] lut_82_select = {
                             in_data[456],
                             in_data[108],
                             in_data[317],
                             in_data[84]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b1100111100001100;
    wire [3:0] lut_83_select = {
                             in_data[291],
                             in_data[258],
                             in_data[613],
                             in_data[320]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b1111000110110000;
    wire [3:0] lut_84_select = {
                             in_data[323],
                             in_data[484],
                             in_data[259],
                             in_data[289]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b0011101100000010;
    wire [3:0] lut_85_select = {
                             in_data[311],
                             in_data[629],
                             in_data[523],
                             in_data[457]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b0011001100110011;
    wire [3:0] lut_86_select = {
                             in_data[469],
                             in_data[496],
                             in_data[335],
                             in_data[333]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b0101010101010101;
    wire [3:0] lut_87_select = {
                             in_data[596],
                             in_data[375],
                             in_data[398],
                             in_data[318]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b1101000011110100;
    wire [3:0] lut_88_select = {
                             in_data[135],
                             in_data[253],
                             in_data[423],
                             in_data[475]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b0000011100010111;
    wire [3:0] lut_89_select = {
                             in_data[283],
                             in_data[117],
                             in_data[265],
                             in_data[623]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1111000010100000;
    wire [3:0] lut_90_select = {
                             in_data[126],
                             in_data[522],
                             in_data[156],
                             in_data[445]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b0111000011110111;
    wire [3:0] lut_91_select = {
                             in_data[200],
                             in_data[406],
                             in_data[194],
                             in_data[468]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1000101110111010;
    wire [3:0] lut_92_select = {
                             in_data[201],
                             in_data[149],
                             in_data[219],
                             in_data[404]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0000111100000101;
    wire [3:0] lut_93_select = {
                             in_data[96],
                             in_data[567],
                             in_data[15],
                             in_data[6]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b0000000011110001;
    wire [3:0] lut_94_select = {
                             in_data[150],
                             in_data[552],
                             in_data[625],
                             in_data[263]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b0011111100100011;
    wire [3:0] lut_95_select = {
                             in_data[85],
                             in_data[458],
                             in_data[542],
                             in_data[553]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b0011001100110011;
    wire [3:0] lut_96_select = {
                             in_data[426],
                             in_data[319],
                             in_data[89],
                             in_data[288]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b0100110111001101;
    wire [3:0] lut_97_select = {
                             in_data[473],
                             in_data[444],
                             in_data[91],
                             in_data[628]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1100010011100100;
    wire [3:0] lut_98_select = {
                             in_data[262],
                             in_data[166],
                             in_data[495],
                             in_data[639]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b0000000011111000;
    wire [3:0] lut_99_select = {
                             in_data[408],
                             in_data[101],
                             in_data[379],
                             in_data[141]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1111000100010001;
    wire [3:0] lut_100_select = {
                             in_data[32],
                             in_data[571],
                             in_data[145],
                             in_data[49]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b0001010000110001;
    wire [3:0] lut_101_select = {
                             in_data[0],
                             in_data[470],
                             in_data[420],
                             in_data[627]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b1010011111100010;
    wire [3:0] lut_102_select = {
                             in_data[213],
                             in_data[393],
                             in_data[86],
                             in_data[142]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1011000011101110;
    wire [3:0] lut_103_select = {
                             in_data[77],
                             in_data[369],
                             in_data[556],
                             in_data[416]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b1110111011101000;
    wire [3:0] lut_104_select = {
                             in_data[622],
                             in_data[314],
                             in_data[237],
                             in_data[356]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1010101011001000;
    wire [3:0] lut_105_select = {
                             in_data[509],
                             in_data[190],
                             in_data[167],
                             in_data[544]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b0000010100010111;
    wire [3:0] lut_106_select = {
                             in_data[578],
                             in_data[340],
                             in_data[462],
                             in_data[427]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b1100000011111100;
    wire [3:0] lut_107_select = {
                             in_data[322],
                             in_data[587],
                             in_data[8],
                             in_data[159]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b0001111100010111;
    wire [3:0] lut_108_select = {
                             in_data[515],
                             in_data[574],
                             in_data[325],
                             in_data[519]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b0000110011001111;
    wire [3:0] lut_109_select = {
                             in_data[436],
                             in_data[125],
                             in_data[593],
                             in_data[29]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b1000100000001110;
    wire [3:0] lut_110_select = {
                             in_data[112],
                             in_data[56],
                             in_data[53],
                             in_data[72]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b1111111100000001;
    wire [3:0] lut_111_select = {
                             in_data[631],
                             in_data[132],
                             in_data[46],
                             in_data[118]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b0010111110111111;
    wire [3:0] lut_112_select = {
                             in_data[243],
                             in_data[216],
                             in_data[276],
                             in_data[206]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b0010001100100010;
    wire [3:0] lut_113_select = {
                             in_data[116],
                             in_data[449],
                             in_data[54],
                             in_data[103]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1100000011010001;
    wire [3:0] lut_114_select = {
                             in_data[610],
                             in_data[14],
                             in_data[361],
                             in_data[274]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b1011101010100000;
    wire [3:0] lut_115_select = {
                             in_data[269],
                             in_data[205],
                             in_data[267],
                             in_data[562]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b0101010101001111;
    wire [3:0] lut_116_select = {
                             in_data[548],
                             in_data[268],
                             in_data[531],
                             in_data[372]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b0000111100001011;
    wire [3:0] lut_117_select = {
                             in_data[499],
                             in_data[225],
                             in_data[634],
                             in_data[67]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1111001010010000;
    wire [3:0] lut_118_select = {
                             in_data[158],
                             in_data[173],
                             in_data[294],
                             in_data[78]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b0001000000110010;
    wire [3:0] lut_119_select = {
                             in_data[328],
                             in_data[421],
                             in_data[527],
                             in_data[90]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b0000000100110101;
    wire [3:0] lut_120_select = {
                             in_data[621],
                             in_data[309],
                             in_data[130],
                             in_data[348]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b1111110111110101;
    wire [3:0] lut_121_select = {
                             in_data[186],
                             in_data[460],
                             in_data[182],
                             in_data[607]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b1011111100000101;
    wire [3:0] lut_122_select = {
                             in_data[566],
                             in_data[48],
                             in_data[308],
                             in_data[241]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b0000001100101111;
    wire [3:0] lut_123_select = {
                             in_data[51],
                             in_data[272],
                             in_data[501],
                             in_data[474]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b1010100011111111;
    wire [3:0] lut_124_select = {
                             in_data[251],
                             in_data[188],
                             in_data[385],
                             in_data[52]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b0000010101011111;
    wire [3:0] lut_125_select = {
                             in_data[636],
                             in_data[535],
                             in_data[2],
                             in_data[195]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b1000000011101110;
    wire [3:0] lut_126_select = {
                             in_data[100],
                             in_data[244],
                             in_data[279],
                             in_data[326]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0011001100110011;
    wire [3:0] lut_127_select = {
                             in_data[177],
                             in_data[18],
                             in_data[355],
                             in_data[597]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b0011011100110011;
    wire [3:0] lut_128_select = {
                             in_data[271],
                             in_data[582],
                             in_data[128],
                             in_data[295]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b0010001000100011;
    wire [3:0] lut_129_select = {
                             in_data[619],
                             in_data[215],
                             in_data[626],
                             in_data[568]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b0000000011101111;
    wire [3:0] lut_130_select = {
                             in_data[57],
                             in_data[378],
                             in_data[329],
                             in_data[347]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b0101110101001101;
    wire [3:0] lut_131_select = {
                             in_data[364],
                             in_data[10],
                             in_data[31],
                             in_data[235]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b0010101100000010;
    wire [3:0] lut_132_select = {
                             in_data[106],
                             in_data[136],
                             in_data[466],
                             in_data[440]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0100010111001111;
    wire [3:0] lut_133_select = {
                             in_data[373],
                             in_data[110],
                             in_data[176],
                             in_data[482]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b1111110011110000;
    wire [3:0] lut_134_select = {
                             in_data[584],
                             in_data[479],
                             in_data[490],
                             in_data[181]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b0001000011110111;
    wire [3:0] lut_135_select = {
                             in_data[485],
                             in_data[559],
                             in_data[428],
                             in_data[102]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b1111111101000000;
    wire [3:0] lut_136_select = {
                             in_data[299],
                             in_data[119],
                             in_data[229],
                             in_data[503]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b1111010011110000;
    wire [3:0] lut_137_select = {
                             in_data[525],
                             in_data[327],
                             in_data[61],
                             in_data[60]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b0100000001010101;
    wire [3:0] lut_138_select = {
                             in_data[76],
                             in_data[511],
                             in_data[534],
                             in_data[75]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b0000010001000101;
    wire [3:0] lut_139_select = {
                             in_data[189],
                             in_data[506],
                             in_data[266],
                             in_data[137]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b1101111111001100;
    wire [3:0] lut_140_select = {
                             in_data[47],
                             in_data[16],
                             in_data[41],
                             in_data[497]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b0111001000000000;
    wire [3:0] lut_141_select = {
                             in_data[236],
                             in_data[601],
                             in_data[303],
                             in_data[443]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b0101011101010101;
    wire [3:0] lut_142_select = {
                             in_data[273],
                             in_data[38],
                             in_data[165],
                             in_data[555]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0000000001001111;
    wire [3:0] lut_143_select = {
                             in_data[611],
                             in_data[592],
                             in_data[304],
                             in_data[352]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b1111001110100000;
    wire [3:0] lut_144_select = {
                             in_data[157],
                             in_data[618],
                             in_data[403],
                             in_data[228]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1100010001000100;
    wire [3:0] lut_145_select = {
                             in_data[44],
                             in_data[3],
                             in_data[405],
                             in_data[387]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1011001011111110;
    wire [3:0] lut_146_select = {
                             in_data[526],
                             in_data[245],
                             in_data[234],
                             in_data[483]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0000000100110011;
    wire [3:0] lut_147_select = {
                             in_data[133],
                             in_data[367],
                             in_data[115],
                             in_data[22]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b1101010111110101;
    wire [3:0] lut_148_select = {
                             in_data[275],
                             in_data[81],
                             in_data[79],
                             in_data[365]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b1111101011111110;
    wire [3:0] lut_149_select = {
                             in_data[417],
                             in_data[353],
                             in_data[134],
                             in_data[174]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b0000010101001111;
    wire [3:0] lut_150_select = {
                             in_data[202],
                             in_data[36],
                             in_data[572],
                             in_data[604]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b1100100011101110;
    wire [3:0] lut_151_select = {
                             in_data[549],
                             in_data[389],
                             in_data[588],
                             in_data[407]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b1011101100110010;
    wire [3:0] lut_152_select = {
                             in_data[489],
                             in_data[576],
                             in_data[540],
                             in_data[297]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1110100011001100;
    wire [3:0] lut_153_select = {
                             in_data[342],
                             in_data[602],
                             in_data[384],
                             in_data[21]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0111000001110001;
    wire [3:0] lut_154_select = {
                             in_data[193],
                             in_data[377],
                             in_data[415],
                             in_data[109]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b1101010111010101;
    wire [3:0] lut_155_select = {
                             in_data[418],
                             in_data[516],
                             in_data[366],
                             in_data[217]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b1111000011111011;
    wire [3:0] lut_156_select = {
                             in_data[620],
                             in_data[399],
                             in_data[435],
                             in_data[305]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b1111111110101010;
    wire [3:0] lut_157_select = {
                             in_data[508],
                             in_data[524],
                             in_data[334],
                             in_data[401]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b1011001011111011;
    wire [3:0] lut_158_select = {
                             in_data[467],
                             in_data[223],
                             in_data[80],
                             in_data[74]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b1010101011101000;
    wire [3:0] lut_159_select = {
                             in_data[33],
                             in_data[73],
                             in_data[363],
                             in_data[306]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b0000111100001111;
    wire [3:0] lut_160_select = {
                             in_data[303],
                             in_data[411],
                             in_data[252],
                             in_data[325]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b0000010000001111;
    wire [3:0] lut_161_select = {
                             in_data[506],
                             in_data[614],
                             in_data[302],
                             in_data[480]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1111011100110001;
    wire [3:0] lut_162_select = {
                             in_data[167],
                             in_data[477],
                             in_data[23],
                             in_data[202]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b0000101000001010;
    wire [3:0] lut_163_select = {
                             in_data[15],
                             in_data[583],
                             in_data[233],
                             in_data[173]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b0101111101001111;
    wire [3:0] lut_164_select = {
                             in_data[565],
                             in_data[331],
                             in_data[538],
                             in_data[487]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b1000110000001100;
    wire [3:0] lut_165_select = {
                             in_data[511],
                             in_data[269],
                             in_data[153],
                             in_data[309]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b1011101010100010;
    wire [3:0] lut_166_select = {
                             in_data[231],
                             in_data[305],
                             in_data[627],
                             in_data[418]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b0010000010111011;
    wire [3:0] lut_167_select = {
                             in_data[621],
                             in_data[120],
                             in_data[208],
                             in_data[488]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b1100110011001100;
    wire [3:0] lut_168_select = {
                             in_data[526],
                             in_data[369],
                             in_data[266],
                             in_data[587]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b1000110000001101;
    wire [3:0] lut_169_select = {
                             in_data[339],
                             in_data[592],
                             in_data[347],
                             in_data[11]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b0101010011111111;
    wire [3:0] lut_170_select = {
                             in_data[373],
                             in_data[527],
                             in_data[612],
                             in_data[358]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b1111101010110010;
    wire [3:0] lut_171_select = {
                             in_data[412],
                             in_data[409],
                             in_data[364],
                             in_data[334]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b0011011101110111;
    wire [3:0] lut_172_select = {
                             in_data[289],
                             in_data[377],
                             in_data[367],
                             in_data[396]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b0010101100100010;
    wire [3:0] lut_173_select = {
                             in_data[333],
                             in_data[384],
                             in_data[152],
                             in_data[122]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b0101111100001101;
    wire [3:0] lut_174_select = {
                             in_data[474],
                             in_data[363],
                             in_data[178],
                             in_data[271]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1001110100001101;
    wire [3:0] lut_175_select = {
                             in_data[43],
                             in_data[539],
                             in_data[124],
                             in_data[256]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b1111011100000000;
    wire [3:0] lut_176_select = {
                             in_data[406],
                             in_data[456],
                             in_data[500],
                             in_data[212]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b1010000011110000;
    wire [3:0] lut_177_select = {
                             in_data[17],
                             in_data[606],
                             in_data[485],
                             in_data[215]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b0111111100000111;
    wire [3:0] lut_178_select = {
                             in_data[564],
                             in_data[216],
                             in_data[442],
                             in_data[435]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b1011000010110011;
    wire [3:0] lut_179_select = {
                             in_data[224],
                             in_data[337],
                             in_data[192],
                             in_data[104]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b1111111100010010;
    wire [3:0] lut_180_select = {
                             in_data[326],
                             in_data[19],
                             in_data[113],
                             in_data[531]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b0101000101010101;
    wire [3:0] lut_181_select = {
                             in_data[290],
                             in_data[187],
                             in_data[566],
                             in_data[35]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b1111000011000000;
    wire [3:0] lut_182_select = {
                             in_data[150],
                             in_data[1],
                             in_data[467],
                             in_data[228]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b0101111101010101;
    wire [3:0] lut_183_select = {
                             in_data[112],
                             in_data[295],
                             in_data[537],
                             in_data[462]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b1000101010001110;
    wire [3:0] lut_184_select = {
                             in_data[610],
                             in_data[482],
                             in_data[628],
                             in_data[620]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b1100010011111100;
    wire [3:0] lut_185_select = {
                             in_data[92],
                             in_data[342],
                             in_data[300],
                             in_data[572]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b1101111111011101;
    wire [3:0] lut_186_select = {
                             in_data[204],
                             in_data[542],
                             in_data[574],
                             in_data[524]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b0100010011011101;
    wire [3:0] lut_187_select = {
                             in_data[26],
                             in_data[513],
                             in_data[308],
                             in_data[503]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b1101010001000000;
    wire [3:0] lut_188_select = {
                             in_data[293],
                             in_data[470],
                             in_data[518],
                             in_data[629]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b0011001100100010;
    wire [3:0] lut_189_select = {
                             in_data[21],
                             in_data[444],
                             in_data[516],
                             in_data[283]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b1111110100000000;
    wire [3:0] lut_190_select = {
                             in_data[454],
                             in_data[354],
                             in_data[179],
                             in_data[407]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b1111100010100000;
    wire [3:0] lut_191_select = {
                             in_data[69],
                             in_data[200],
                             in_data[545],
                             in_data[590]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b1111110100010000;
    wire [3:0] lut_192_select = {
                             in_data[162],
                             in_data[429],
                             in_data[630],
                             in_data[54]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b0100000011111100;
    wire [3:0] lut_193_select = {
                             in_data[371],
                             in_data[346],
                             in_data[195],
                             in_data[370]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0100000101010001;
    wire [3:0] lut_194_select = {
                             in_data[169],
                             in_data[552],
                             in_data[25],
                             in_data[199]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b1111010101010001;
    wire [3:0] lut_195_select = {
                             in_data[413],
                             in_data[157],
                             in_data[495],
                             in_data[555]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b1111011101010001;
    wire [3:0] lut_196_select = {
                             in_data[341],
                             in_data[196],
                             in_data[458],
                             in_data[359]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b0000000000111110;
    wire [3:0] lut_197_select = {
                             in_data[558],
                             in_data[595],
                             in_data[97],
                             in_data[395]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b1100100011001110;
    wire [3:0] lut_198_select = {
                             in_data[240],
                             in_data[291],
                             in_data[568],
                             in_data[533]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b0000000010001111;
    wire [3:0] lut_199_select = {
                             in_data[48],
                             in_data[41],
                             in_data[553],
                             in_data[222]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b1010101011111111;
    wire [3:0] lut_200_select = {
                             in_data[338],
                             in_data[351],
                             in_data[391],
                             in_data[129]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b0100010011000100;
    wire [3:0] lut_201_select = {
                             in_data[519],
                             in_data[479],
                             in_data[306],
                             in_data[138]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b1011001000100000;
    wire [3:0] lut_202_select = {
                             in_data[447],
                             in_data[414],
                             in_data[160],
                             in_data[284]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b1100000011000000;
    wire [3:0] lut_203_select = {
                             in_data[180],
                             in_data[286],
                             in_data[489],
                             in_data[76]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b0000000000001100;
    wire [3:0] lut_204_select = {
                             in_data[64],
                             in_data[163],
                             in_data[410],
                             in_data[101]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b0011001100110011;
    wire [3:0] lut_205_select = {
                             in_data[312],
                             in_data[445],
                             in_data[426],
                             in_data[637]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b1010001010100000;
    wire [3:0] lut_206_select = {
                             in_data[143],
                             in_data[625],
                             in_data[455],
                             in_data[151]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b1111010000000000;
    wire [3:0] lut_207_select = {
                             in_data[144],
                             in_data[175],
                             in_data[415],
                             in_data[299]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1110101011101000;
    wire [3:0] lut_208_select = {
                             in_data[203],
                             in_data[55],
                             in_data[402],
                             in_data[603]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b0011011101110111;
    wire [3:0] lut_209_select = {
                             in_data[509],
                             in_data[2],
                             in_data[382],
                             in_data[248]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b1000101000001010;
    wire [3:0] lut_210_select = {
                             in_data[322],
                             in_data[438],
                             in_data[83],
                             in_data[514]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b0010001110111111;
    wire [3:0] lut_211_select = {
                             in_data[457],
                             in_data[490],
                             in_data[66],
                             in_data[381]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b0011111100001011;
    wire [3:0] lut_212_select = {
                             in_data[185],
                             in_data[401],
                             in_data[298],
                             in_data[99]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b1100010011111101;
    wire [3:0] lut_213_select = {
                             in_data[237],
                             in_data[265],
                             in_data[98],
                             in_data[523]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1011001110110010;
    wire [3:0] lut_214_select = {
                             in_data[344],
                             in_data[602],
                             in_data[343],
                             in_data[235]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b1011101100100010;
    wire [3:0] lut_215_select = {
                             in_data[548],
                             in_data[605],
                             in_data[349],
                             in_data[634]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b1101110101011101;
    wire [3:0] lut_216_select = {
                             in_data[465],
                             in_data[130],
                             in_data[255],
                             in_data[89]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b1111101000000010;
    wire [3:0] lut_217_select = {
                             in_data[471],
                             in_data[596],
                             in_data[194],
                             in_data[582]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b1010000010111011;
    wire [3:0] lut_218_select = {
                             in_data[218],
                             in_data[90],
                             in_data[608],
                             in_data[588]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b0011011100000011;
    wire [3:0] lut_219_select = {
                             in_data[374],
                             in_data[546],
                             in_data[205],
                             in_data[51]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b0010101110101011;
    wire [3:0] lut_220_select = {
                             in_data[77],
                             in_data[601],
                             in_data[521],
                             in_data[5]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b0111111100000111;
    wire [3:0] lut_221_select = {
                             in_data[8],
                             in_data[310],
                             in_data[247],
                             in_data[464]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b0000100010111111;
    wire [3:0] lut_222_select = {
                             in_data[615],
                             in_data[221],
                             in_data[109],
                             in_data[183]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1000111111001100;
    wire [3:0] lut_223_select = {
                             in_data[146],
                             in_data[107],
                             in_data[356],
                             in_data[174]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b1000111010001000;
    wire [3:0] lut_224_select = {
                             in_data[379],
                             in_data[619],
                             in_data[313],
                             in_data[376]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b1110111110101010;
    wire [3:0] lut_225_select = {
                             in_data[188],
                             in_data[473],
                             in_data[557],
                             in_data[281]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1111101111000000;
    wire [3:0] lut_226_select = {
                             in_data[9],
                             in_data[393],
                             in_data[505],
                             in_data[176]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b0000101111111111;
    wire [3:0] lut_227_select = {
                             in_data[534],
                             in_data[448],
                             in_data[133],
                             in_data[139]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b1010101011111111;
    wire [3:0] lut_228_select = {
                             in_data[361],
                             in_data[206],
                             in_data[626],
                             in_data[241]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b1100010011101110;
    wire [3:0] lut_229_select = {
                             in_data[123],
                             in_data[633],
                             in_data[128],
                             in_data[125]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b0010000011110010;
    wire [3:0] lut_230_select = {
                             in_data[554],
                             in_data[436],
                             in_data[14],
                             in_data[148]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b1000100010101110;
    wire [3:0] lut_231_select = {
                             in_data[400],
                             in_data[451],
                             in_data[589],
                             in_data[323]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b1100111100001101;
    wire [3:0] lut_232_select = {
                             in_data[461],
                             in_data[168],
                             in_data[74],
                             in_data[106]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b0000000001011100;
    wire [3:0] lut_233_select = {
                             in_data[385],
                             in_data[282],
                             in_data[632],
                             in_data[0]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b1010100010110000;
    wire [3:0] lut_234_select = {
                             in_data[262],
                             in_data[257],
                             in_data[280],
                             in_data[186]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b1110100011111110;
    wire [3:0] lut_235_select = {
                             in_data[198],
                             in_data[631],
                             in_data[484],
                             in_data[131]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b0010101000000010;
    wire [3:0] lut_236_select = {
                             in_data[60],
                             in_data[498],
                             in_data[304],
                             in_data[551]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b1110101000001000;
    wire [3:0] lut_237_select = {
                             in_data[108],
                             in_data[159],
                             in_data[12],
                             in_data[201]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b1010111100001011;
    wire [3:0] lut_238_select = {
                             in_data[317],
                             in_data[18],
                             in_data[556],
                             in_data[115]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0111011101110001;
    wire [3:0] lut_239_select = {
                             in_data[145],
                             in_data[586],
                             in_data[604],
                             in_data[316]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b1110100011110011;
    wire [3:0] lut_240_select = {
                             in_data[86],
                             in_data[190],
                             in_data[261],
                             in_data[184]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b0101000011110000;
    wire [3:0] lut_241_select = {
                             in_data[57],
                             in_data[264],
                             in_data[353],
                             in_data[622]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b0011000010110000;
    wire [3:0] lut_242_select = {
                             in_data[31],
                             in_data[4],
                             in_data[37],
                             in_data[177]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b1000000010101000;
    wire [3:0] lut_243_select = {
                             in_data[549],
                             in_data[397],
                             in_data[268],
                             in_data[242]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b1111111011101010;
    wire [3:0] lut_244_select = {
                             in_data[501],
                             in_data[78],
                             in_data[253],
                             in_data[81]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b0101001100110001;
    wire [3:0] lut_245_select = {
                             in_data[100],
                             in_data[191],
                             in_data[217],
                             in_data[386]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b1101110101001100;
    wire [3:0] lut_246_select = {
                             in_data[529],
                             in_data[102],
                             in_data[504],
                             in_data[563]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b0011001101110001;
    wire [3:0] lut_247_select = {
                             in_data[497],
                             in_data[278],
                             in_data[91],
                             in_data[223]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b0101000001010001;
    wire [3:0] lut_248_select = {
                             in_data[434],
                             in_data[33],
                             in_data[611],
                             in_data[46]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b0011001100111111;
    wire [3:0] lut_249_select = {
                             in_data[535],
                             in_data[577],
                             in_data[493],
                             in_data[126]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b1111100011111110;
    wire [3:0] lut_250_select = {
                             in_data[491],
                             in_data[79],
                             in_data[36],
                             in_data[460]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b0011101110111011;
    wire [3:0] lut_251_select = {
                             in_data[547],
                             in_data[450],
                             in_data[517],
                             in_data[210]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b0101000101010001;
    wire [3:0] lut_252_select = {
                             in_data[387],
                             in_data[49],
                             in_data[431],
                             in_data[638]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b0000110001111111;
    wire [3:0] lut_253_select = {
                             in_data[425],
                             in_data[368],
                             in_data[296],
                             in_data[567]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b1011111000101110;
    wire [3:0] lut_254_select = {
                             in_data[439],
                             in_data[238],
                             in_data[29],
                             in_data[392]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b1100110011001101;
    wire [3:0] lut_255_select = {
                             in_data[475],
                             in_data[335],
                             in_data[559],
                             in_data[249]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b0101010100010111;
    wire [3:0] lut_256_select = {
                             in_data[576],
                             in_data[52],
                             in_data[544],
                             in_data[61]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b0000111100000100;
    wire [3:0] lut_257_select = {
                             in_data[319],
                             in_data[117],
                             in_data[16],
                             in_data[272]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b1111000011111111;
    wire [3:0] lut_258_select = {
                             in_data[70],
                             in_data[225],
                             in_data[32],
                             in_data[609]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b1111001011111011;
    wire [3:0] lut_259_select = {
                             in_data[562],
                             in_data[580],
                             in_data[383],
                             in_data[42]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b0101011101000101;
    wire [3:0] lut_260_select = {
                             in_data[95],
                             in_data[593],
                             in_data[259],
                             in_data[616]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b0010101000101011;
    wire [3:0] lut_261_select = {
                             in_data[75],
                             in_data[147],
                             in_data[449],
                             in_data[599]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b1111000011111111;
    wire [3:0] lut_262_select = {
                             in_data[244],
                             in_data[229],
                             in_data[132],
                             in_data[294]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b0111000101110111;
    wire [3:0] lut_263_select = {
                             in_data[348],
                             in_data[598],
                             in_data[230],
                             in_data[571]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b1111000000110010;
    wire [3:0] lut_264_select = {
                             in_data[7],
                             in_data[543],
                             in_data[419],
                             in_data[466]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b0001101100000010;
    wire [3:0] lut_265_select = {
                             in_data[440],
                             in_data[352],
                             in_data[22],
                             in_data[20]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1111010101010000;
    wire [3:0] lut_266_select = {
                             in_data[260],
                             in_data[245],
                             in_data[607],
                             in_data[428]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b1011101011111011;
    wire [3:0] lut_267_select = {
                             in_data[236],
                             in_data[578],
                             in_data[137],
                             in_data[416]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1110000011111100;
    wire [3:0] lut_268_select = {
                             in_data[591],
                             in_data[581],
                             in_data[618],
                             in_data[82]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0111011101010101;
    wire [3:0] lut_269_select = {
                             in_data[536],
                             in_data[88],
                             in_data[105],
                             in_data[579]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b1100100011001000;
    wire [3:0] lut_270_select = {
                             in_data[408],
                             in_data[127],
                             in_data[452],
                             in_data[389]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b1011101100110011;
    wire [3:0] lut_271_select = {
                             in_data[314],
                             in_data[424],
                             in_data[510],
                             in_data[525]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b1111010111110101;
    wire [3:0] lut_272_select = {
                             in_data[315],
                             in_data[404],
                             in_data[24],
                             in_data[372]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b1010111100001010;
    wire [3:0] lut_273_select = {
                             in_data[350],
                             in_data[327],
                             in_data[446],
                             in_data[10]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b0100111101001101;
    wire [3:0] lut_274_select = {
                             in_data[30],
                             in_data[623],
                             in_data[85],
                             in_data[496]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b0010101000100010;
    wire [3:0] lut_275_select = {
                             in_data[380],
                             in_data[332],
                             in_data[492],
                             in_data[297]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b1111000101000000;
    wire [3:0] lut_276_select = {
                             in_data[254],
                             in_data[246],
                             in_data[63],
                             in_data[617]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b1111110111001100;
    wire [3:0] lut_277_select = {
                             in_data[39],
                             in_data[324],
                             in_data[53],
                             in_data[94]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b1000110010001000;
    wire [3:0] lut_278_select = {
                             in_data[430],
                             in_data[219],
                             in_data[378],
                             in_data[243]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b0101010101010100;
    wire [3:0] lut_279_select = {
                             in_data[357],
                             in_data[321],
                             in_data[267],
                             in_data[522]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b1101010111010100;
    wire [3:0] lut_280_select = {
                             in_data[181],
                             in_data[156],
                             in_data[486],
                             in_data[398]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b1010111000001000;
    wire [3:0] lut_281_select = {
                             in_data[158],
                             in_data[481],
                             in_data[80],
                             in_data[44]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b0000110111111111;
    wire [3:0] lut_282_select = {
                             in_data[67],
                             in_data[232],
                             in_data[171],
                             in_data[189]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b1110100010100000;
    wire [3:0] lut_283_select = {
                             in_data[561],
                             in_data[530],
                             in_data[441],
                             in_data[275]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b0000010011001101;
    wire [3:0] lut_284_select = {
                             in_data[65],
                             in_data[427],
                             in_data[585],
                             in_data[355]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b0010111100001011;
    wire [3:0] lut_285_select = {
                             in_data[512],
                             in_data[165],
                             in_data[140],
                             in_data[6]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b1110111011101110;
    wire [3:0] lut_286_select = {
                             in_data[258],
                             in_data[154],
                             in_data[285],
                             in_data[111]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b1100000011010000;
    wire [3:0] lut_287_select = {
                             in_data[520],
                             in_data[72],
                             in_data[155],
                             in_data[320]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b0110010001111111;
    wire [3:0] lut_288_select = {
                             in_data[116],
                             in_data[277],
                             in_data[502],
                             in_data[273]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b1110111010101000;
    wire [3:0] lut_289_select = {
                             in_data[211],
                             in_data[453],
                             in_data[68],
                             in_data[28]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b0111011100000001;
    wire [3:0] lut_290_select = {
                             in_data[110],
                             in_data[234],
                             in_data[172],
                             in_data[213]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b1000110110001110;
    wire [3:0] lut_291_select = {
                             in_data[170],
                             in_data[56],
                             in_data[494],
                             in_data[399]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b0000111100001111;
    wire [3:0] lut_292_select = {
                             in_data[600],
                             in_data[311],
                             in_data[443],
                             in_data[47]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b1011101010101010;
    wire [3:0] lut_293_select = {
                             in_data[214],
                             in_data[38],
                             in_data[636],
                             in_data[345]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1011111100000010;
    wire [3:0] lut_294_select = {
                             in_data[118],
                             in_data[274],
                             in_data[478],
                             in_data[250]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b0111000101110111;
    wire [3:0] lut_295_select = {
                             in_data[469],
                             in_data[119],
                             in_data[483],
                             in_data[197]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b1100000011111100;
    wire [3:0] lut_296_select = {
                             in_data[71],
                             in_data[135],
                             in_data[394],
                             in_data[182]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b1110111100001100;
    wire [3:0] lut_297_select = {
                             in_data[330],
                             in_data[575],
                             in_data[507],
                             in_data[239]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b0011001000100000;
    wire [3:0] lut_298_select = {
                             in_data[73],
                             in_data[329],
                             in_data[149],
                             in_data[422]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b1111100011110000;
    wire [3:0] lut_299_select = {
                             in_data[573],
                             in_data[276],
                             in_data[433],
                             in_data[624]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b1010001010101010;
    wire [3:0] lut_300_select = {
                             in_data[437],
                             in_data[594],
                             in_data[468],
                             in_data[263]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b1010001010110011;
    wire [3:0] lut_301_select = {
                             in_data[360],
                             in_data[220],
                             in_data[142],
                             in_data[318]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b1111110011001000;
    wire [3:0] lut_302_select = {
                             in_data[540],
                             in_data[432],
                             in_data[62],
                             in_data[34]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b1010111110101111;
    wire [3:0] lut_303_select = {
                             in_data[417],
                             in_data[365],
                             in_data[459],
                             in_data[528]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b0100111100010111;
    wire [3:0] lut_304_select = {
                             in_data[45],
                             in_data[532],
                             in_data[164],
                             in_data[50]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b1111000011111000;
    wire [3:0] lut_305_select = {
                             in_data[307],
                             in_data[301],
                             in_data[114],
                             in_data[93]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b0100110001000100;
    wire [3:0] lut_306_select = {
                             in_data[423],
                             in_data[166],
                             in_data[388],
                             in_data[27]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b0000000110111111;
    wire [3:0] lut_307_select = {
                             in_data[84],
                             in_data[40],
                             in_data[403],
                             in_data[59]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b0000010101010101;
    wire [3:0] lut_308_select = {
                             in_data[96],
                             in_data[463],
                             in_data[476],
                             in_data[209]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b0000010101000100;
    wire [3:0] lut_309_select = {
                             in_data[635],
                             in_data[508],
                             in_data[639],
                             in_data[193]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b0000000011000000;
    wire [3:0] lut_310_select = {
                             in_data[134],
                             in_data[103],
                             in_data[226],
                             in_data[613]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b0101010101000000;
    wire [3:0] lut_311_select = {
                             in_data[121],
                             in_data[270],
                             in_data[570],
                             in_data[13]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1110111100001111;
    wire [3:0] lut_312_select = {
                             in_data[161],
                             in_data[3],
                             in_data[328],
                             in_data[288]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b0101000111110000;
    wire [3:0] lut_313_select = {
                             in_data[499],
                             in_data[141],
                             in_data[362],
                             in_data[227]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b1010101000001000;
    wire [3:0] lut_314_select = {
                             in_data[472],
                             in_data[560],
                             in_data[550],
                             in_data[136]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b1010100010101000;
    wire [3:0] lut_315_select = {
                             in_data[597],
                             in_data[287],
                             in_data[279],
                             in_data[569]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b0000000010101011;
    wire [3:0] lut_316_select = {
                             in_data[366],
                             in_data[336],
                             in_data[541],
                             in_data[420]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b1111000010110000;
    wire [3:0] lut_317_select = {
                             in_data[405],
                             in_data[515],
                             in_data[292],
                             in_data[584]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0000000000001111;
    wire [3:0] lut_318_select = {
                             in_data[87],
                             in_data[58],
                             in_data[421],
                             in_data[340]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b0001001101111111;
    wire [3:0] lut_319_select = {
                             in_data[375],
                             in_data[207],
                             in_data[251],
                             in_data[390]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b0111011100110001;
    wire [3:0] lut_320_select = {
                             in_data[615],
                             in_data[366],
                             in_data[52],
                             in_data[235]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0100010101001101;
    wire [3:0] lut_321_select = {
                             in_data[477],
                             in_data[561],
                             in_data[273],
                             in_data[291]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b1100000011111111;
    wire [3:0] lut_322_select = {
                             in_data[468],
                             in_data[338],
                             in_data[219],
                             in_data[451]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b1111000100000000;
    wire [3:0] lut_323_select = {
                             in_data[70],
                             in_data[398],
                             in_data[414],
                             in_data[147]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b1000111000000000;
    wire [3:0] lut_324_select = {
                             in_data[552],
                             in_data[153],
                             in_data[631],
                             in_data[108]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b0000101000001111;
    wire [3:0] lut_325_select = {
                             in_data[349],
                             in_data[433],
                             in_data[154],
                             in_data[324]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b1111010011010100;
    wire [3:0] lut_326_select = {
                             in_data[55],
                             in_data[21],
                             in_data[590],
                             in_data[353]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b0000000010111011;
    wire [3:0] lut_327_select = {
                             in_data[286],
                             in_data[604],
                             in_data[464],
                             in_data[405]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b0111111101110000;
    wire [3:0] lut_328_select = {
                             in_data[429],
                             in_data[35],
                             in_data[133],
                             in_data[438]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b0000010100010101;
    wire [3:0] lut_329_select = {
                             in_data[471],
                             in_data[166],
                             in_data[305],
                             in_data[387]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b1111100011101000;
    wire [3:0] lut_330_select = {
                             in_data[453],
                             in_data[634],
                             in_data[90],
                             in_data[8]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b0000000100000011;
    wire [3:0] lut_331_select = {
                             in_data[180],
                             in_data[268],
                             in_data[174],
                             in_data[51]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b1110111010101010;
    wire [3:0] lut_332_select = {
                             in_data[53],
                             in_data[261],
                             in_data[298],
                             in_data[56]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b1111111100001010;
    wire [3:0] lut_333_select = {
                             in_data[524],
                             in_data[170],
                             in_data[132],
                             in_data[284]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b1000110011001110;
    wire [3:0] lut_334_select = {
                             in_data[421],
                             in_data[584],
                             in_data[345],
                             in_data[500]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0010101100101011;
    wire [3:0] lut_335_select = {
                             in_data[136],
                             in_data[206],
                             in_data[44],
                             in_data[274]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b1111101110101000;
    wire [3:0] lut_336_select = {
                             in_data[550],
                             in_data[517],
                             in_data[49],
                             in_data[583]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b1010101000101010;
    wire [3:0] lut_337_select = {
                             in_data[97],
                             in_data[603],
                             in_data[490],
                             in_data[367]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b0000010100000101;
    wire [3:0] lut_338_select = {
                             in_data[62],
                             in_data[492],
                             in_data[466],
                             in_data[611]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b1010101010101010;
    wire [3:0] lut_339_select = {
                             in_data[616],
                             in_data[225],
                             in_data[446],
                             in_data[276]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b1111000111110100;
    wire [3:0] lut_340_select = {
                             in_data[80],
                             in_data[407],
                             in_data[502],
                             in_data[327]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b1010111000001000;
    wire [3:0] lut_341_select = {
                             in_data[242],
                             in_data[119],
                             in_data[110],
                             in_data[222]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b1011001010100000;
    wire [3:0] lut_342_select = {
                             in_data[486],
                             in_data[200],
                             in_data[636],
                             in_data[272]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b0100111000001110;
    wire [3:0] lut_343_select = {
                             in_data[211],
                             in_data[168],
                             in_data[411],
                             in_data[114]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1010000010100000;
    wire [3:0] lut_344_select = {
                             in_data[428],
                             in_data[511],
                             in_data[248],
                             in_data[107]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b0100111100101111;
    wire [3:0] lut_345_select = {
                             in_data[176],
                             in_data[165],
                             in_data[295],
                             in_data[385]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b1000100011111111;
    wire [3:0] lut_346_select = {
                             in_data[104],
                             in_data[263],
                             in_data[410],
                             in_data[0]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b1100110011001110;
    wire [3:0] lut_347_select = {
                             in_data[621],
                             in_data[565],
                             in_data[279],
                             in_data[356]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0000000100010111;
    wire [3:0] lut_348_select = {
                             in_data[193],
                             in_data[521],
                             in_data[149],
                             in_data[11]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b0010111101111111;
    wire [3:0] lut_349_select = {
                             in_data[232],
                             in_data[607],
                             in_data[637],
                             in_data[573]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b0111001101110001;
    wire [3:0] lut_350_select = {
                             in_data[626],
                             in_data[37],
                             in_data[638],
                             in_data[60]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b1111110000000000;
    wire [3:0] lut_351_select = {
                             in_data[150],
                             in_data[197],
                             in_data[533],
                             in_data[333]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b0111011101110101;
    wire [3:0] lut_352_select = {
                             in_data[258],
                             in_data[39],
                             in_data[138],
                             in_data[98]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b1111001100110000;
    wire [3:0] lut_353_select = {
                             in_data[31],
                             in_data[280],
                             in_data[470],
                             in_data[74]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b0000001001111111;
    wire [3:0] lut_354_select = {
                             in_data[59],
                             in_data[518],
                             in_data[192],
                             in_data[159]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b0000101011111111;
    wire [3:0] lut_355_select = {
                             in_data[337],
                             in_data[188],
                             in_data[121],
                             in_data[409]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b0101000101110000;
    wire [3:0] lut_356_select = {
                             in_data[122],
                             in_data[5],
                             in_data[13],
                             in_data[294]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b0010101100100010;
    wire [3:0] lut_357_select = {
                             in_data[113],
                             in_data[506],
                             in_data[134],
                             in_data[450]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b0100111100010111;
    wire [3:0] lut_358_select = {
                             in_data[162],
                             in_data[539],
                             in_data[260],
                             in_data[443]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b0000101000000111;
    wire [3:0] lut_359_select = {
                             in_data[633],
                             in_data[448],
                             in_data[553],
                             in_data[283]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b1000000011000000;
    wire [3:0] lut_360_select = {
                             in_data[36],
                             in_data[529],
                             in_data[83],
                             in_data[308]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b0111111100000111;
    wire [3:0] lut_361_select = {
                             in_data[190],
                             in_data[544],
                             in_data[579],
                             in_data[434]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b0100111000001000;
    wire [3:0] lut_362_select = {
                             in_data[16],
                             in_data[538],
                             in_data[447],
                             in_data[473]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b0001111101110111;
    wire [3:0] lut_363_select = {
                             in_data[632],
                             in_data[559],
                             in_data[230],
                             in_data[396]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b0001111101011111;
    wire [3:0] lut_364_select = {
                             in_data[600],
                             in_data[493],
                             in_data[487],
                             in_data[424]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b1100110011001100;
    wire [3:0] lut_365_select = {
                             in_data[478],
                             in_data[588],
                             in_data[381],
                             in_data[129]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b0101010101110000;
    wire [3:0] lut_366_select = {
                             in_data[370],
                             in_data[25],
                             in_data[629],
                             in_data[292]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b1110111010101110;
    wire [3:0] lut_367_select = {
                             in_data[93],
                             in_data[256],
                             in_data[560],
                             in_data[392]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b1111110111101110;
    wire [3:0] lut_368_select = {
                             in_data[509],
                             in_data[397],
                             in_data[460],
                             in_data[40]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b0000000011111111;
    wire [3:0] lut_369_select = {
                             in_data[505],
                             in_data[599],
                             in_data[557],
                             in_data[362]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b1011100010100000;
    wire [3:0] lut_370_select = {
                             in_data[281],
                             in_data[365],
                             in_data[204],
                             in_data[311]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b1110100011001000;
    wire [3:0] lut_371_select = {
                             in_data[580],
                             in_data[540],
                             in_data[419],
                             in_data[507]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b1101010001110101;
    wire [3:0] lut_372_select = {
                             in_data[253],
                             in_data[306],
                             in_data[569],
                             in_data[556]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b0000111111011111;
    wire [3:0] lut_373_select = {
                             in_data[564],
                             in_data[151],
                             in_data[304],
                             in_data[426]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b1011001110110011;
    wire [3:0] lut_374_select = {
                             in_data[47],
                             in_data[329],
                             in_data[30],
                             in_data[578]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b0101000001010101;
    wire [3:0] lut_375_select = {
                             in_data[610],
                             in_data[591],
                             in_data[6],
                             in_data[315]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b1000110011001110;
    wire [3:0] lut_376_select = {
                             in_data[501],
                             in_data[290],
                             in_data[627],
                             in_data[449]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b0101111100001111;
    wire [3:0] lut_377_select = {
                             in_data[562],
                             in_data[71],
                             in_data[437],
                             in_data[313]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b0101110101011101;
    wire [3:0] lut_378_select = {
                             in_data[618],
                             in_data[476],
                             in_data[91],
                             in_data[140]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1111110011001100;
    wire [3:0] lut_379_select = {
                             in_data[465],
                             in_data[251],
                             in_data[628],
                             in_data[322]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b0100010001010101;
    wire [3:0] lut_380_select = {
                             in_data[625],
                             in_data[339],
                             in_data[452],
                             in_data[459]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b0100000011001100;
    wire [3:0] lut_381_select = {
                             in_data[217],
                             in_data[455],
                             in_data[250],
                             in_data[14]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b0000000011111111;
    wire [3:0] lut_382_select = {
                             in_data[359],
                             in_data[467],
                             in_data[67],
                             in_data[307]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b0011101100100011;
    wire [3:0] lut_383_select = {
                             in_data[495],
                             in_data[109],
                             in_data[207],
                             in_data[555]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0100010111001101;
    wire [3:0] lut_384_select = {
                             in_data[297],
                             in_data[328],
                             in_data[360],
                             in_data[194]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b1111111110001000;
    wire [3:0] lut_385_select = {
                             in_data[474],
                             in_data[24],
                             in_data[208],
                             in_data[128]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b0000000011110000;
    wire [3:0] lut_386_select = {
                             in_data[257],
                             in_data[143],
                             in_data[382],
                             in_data[456]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b1101110111001100;
    wire [3:0] lut_387_select = {
                             in_data[420],
                             in_data[185],
                             in_data[227],
                             in_data[617]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b0001000100110011;
    wire [3:0] lut_388_select = {
                             in_data[177],
                             in_data[534],
                             in_data[285],
                             in_data[318]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b1100110101000100;
    wire [3:0] lut_389_select = {
                             in_data[479],
                             in_data[175],
                             in_data[369],
                             in_data[54]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b1010101010001010;
    wire [3:0] lut_390_select = {
                             in_data[43],
                             in_data[519],
                             in_data[388],
                             in_data[34]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b0001000100010111;
    wire [3:0] lut_391_select = {
                             in_data[2],
                             in_data[301],
                             in_data[224],
                             in_data[567]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b0010101000100010;
    wire [3:0] lut_392_select = {
                             in_data[440],
                             in_data[247],
                             in_data[220],
                             in_data[148]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b1110101010101010;
    wire [3:0] lut_393_select = {
                             in_data[82],
                             in_data[117],
                             in_data[77],
                             in_data[179]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b1010111100101111;
    wire [3:0] lut_394_select = {
                             in_data[264],
                             in_data[321],
                             in_data[46],
                             in_data[233]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b1110101010001000;
    wire [3:0] lut_395_select = {
                             in_data[214],
                             in_data[12],
                             in_data[347],
                             in_data[103]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b1100111000001110;
    wire [3:0] lut_396_select = {
                             in_data[244],
                             in_data[296],
                             in_data[497],
                             in_data[619]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b0000110000001100;
    wire [3:0] lut_397_select = {
                             in_data[542],
                             in_data[606],
                             in_data[293],
                             in_data[520]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b1111000011111010;
    wire [3:0] lut_398_select = {
                             in_data[575],
                             in_data[605],
                             in_data[65],
                             in_data[287]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b0101011100000101;
    wire [3:0] lut_399_select = {
                             in_data[394],
                             in_data[601],
                             in_data[335],
                             in_data[445]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b1011101000000000;
    wire [3:0] lut_400_select = {
                             in_data[237],
                             in_data[203],
                             in_data[212],
                             in_data[302]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b0011001100010011;
    wire [3:0] lut_401_select = {
                             in_data[255],
                             in_data[88],
                             in_data[23],
                             in_data[422]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b1100110011001100;
    wire [3:0] lut_402_select = {
                             in_data[401],
                             in_data[68],
                             in_data[7],
                             in_data[81]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b0000010100001101;
    wire [3:0] lut_403_select = {
                             in_data[418],
                             in_data[95],
                             in_data[341],
                             in_data[130]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b1011001011110000;
    wire [3:0] lut_404_select = {
                             in_data[271],
                             in_data[288],
                             in_data[19],
                             in_data[123]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b1100110011111101;
    wire [3:0] lut_405_select = {
                             in_data[489],
                             in_data[131],
                             in_data[442],
                             in_data[549]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0101000101010101;
    wire [3:0] lut_406_select = {
                             in_data[229],
                             in_data[375],
                             in_data[379],
                             in_data[576]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b0000010101010101;
    wire [3:0] lut_407_select = {
                             in_data[558],
                             in_data[323],
                             in_data[213],
                             in_data[20]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b1100000011000000;
    wire [3:0] lut_408_select = {
                             in_data[9],
                             in_data[581],
                             in_data[320],
                             in_data[196]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b0000000000001111;
    wire [3:0] lut_409_select = {
                             in_data[157],
                             in_data[566],
                             in_data[231],
                             in_data[309]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b0000000010101111;
    wire [3:0] lut_410_select = {
                             in_data[319],
                             in_data[238],
                             in_data[28],
                             in_data[386]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b1100000011101000;
    wire [3:0] lut_411_select = {
                             in_data[523],
                             in_data[639],
                             in_data[202],
                             in_data[331]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b0001011101111111;
    wire [3:0] lut_412_select = {
                             in_data[522],
                             in_data[312],
                             in_data[350],
                             in_data[73]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b1100110011101110;
    wire [3:0] lut_413_select = {
                             in_data[585],
                             in_data[326],
                             in_data[535],
                             in_data[571]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0001000011110111;
    wire [3:0] lut_414_select = {
                             in_data[594],
                             in_data[205],
                             in_data[514],
                             in_data[317]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b1111001111110011;
    wire [3:0] lut_415_select = {
                             in_data[289],
                             in_data[547],
                             in_data[105],
                             in_data[589]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b1101110111111111;
    wire [3:0] lut_416_select = {
                             in_data[416],
                             in_data[184],
                             in_data[115],
                             in_data[45]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b1100111010101110;
    wire [3:0] lut_417_select = {
                             in_data[310],
                             in_data[76],
                             in_data[223],
                             in_data[336]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b0000000011110101;
    wire [3:0] lut_418_select = {
                             in_data[259],
                             in_data[361],
                             in_data[15],
                             in_data[602]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b1111001110110000;
    wire [3:0] lut_419_select = {
                             in_data[403],
                             in_data[475],
                             in_data[404],
                             in_data[92]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b1100111000001000;
    wire [3:0] lut_420_select = {
                             in_data[596],
                             in_data[270],
                             in_data[161],
                             in_data[332]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b0000000000110011;
    wire [3:0] lut_421_select = {
                             in_data[498],
                             in_data[541],
                             in_data[512],
                             in_data[572]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b1100110011000000;
    wire [3:0] lut_422_select = {
                             in_data[254],
                             in_data[526],
                             in_data[84],
                             in_data[357]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b1110100011101100;
    wire [3:0] lut_423_select = {
                             in_data[152],
                             in_data[482],
                             in_data[463],
                             in_data[574]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b0010100000101011;
    wire [3:0] lut_424_select = {
                             in_data[496],
                             in_data[156],
                             in_data[169],
                             in_data[430]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b0001000001010001;
    wire [3:0] lut_425_select = {
                             in_data[377],
                             in_data[348],
                             in_data[432],
                             in_data[218]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b0000011100000011;
    wire [3:0] lut_426_select = {
                             in_data[537],
                             in_data[142],
                             in_data[358],
                             in_data[112]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b0010101010101011;
    wire [3:0] lut_427_select = {
                             in_data[503],
                             in_data[485],
                             in_data[29],
                             in_data[536]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b0111011100100101;
    wire [3:0] lut_428_select = {
                             in_data[508],
                             in_data[346],
                             in_data[491],
                             in_data[368]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b1000111011101111;
    wire [3:0] lut_429_select = {
                             in_data[425],
                             in_data[191],
                             in_data[245],
                             in_data[144]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b0010101110111111;
    wire [3:0] lut_430_select = {
                             in_data[620],
                             in_data[554],
                             in_data[515],
                             in_data[163]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b0000000011111111;
    wire [3:0] lut_431_select = {
                             in_data[125],
                             in_data[635],
                             in_data[278],
                             in_data[395]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b0111000101110011;
    wire [3:0] lut_432_select = {
                             in_data[171],
                             in_data[436],
                             in_data[390],
                             in_data[355]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b1110111111001110;
    wire [3:0] lut_433_select = {
                             in_data[528],
                             in_data[444],
                             in_data[137],
                             in_data[316]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b1111100011111101;
    wire [3:0] lut_434_select = {
                             in_data[372],
                             in_data[38],
                             in_data[187],
                             in_data[141]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b1011101010101000;
    wire [3:0] lut_435_select = {
                             in_data[622],
                             in_data[85],
                             in_data[300],
                             in_data[234]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b0011000100110001;
    wire [3:0] lut_436_select = {
                             in_data[344],
                             in_data[215],
                             in_data[488],
                             in_data[408]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b0000011100011111;
    wire [3:0] lut_437_select = {
                             in_data[595],
                             in_data[94],
                             in_data[181],
                             in_data[461]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b0001000001110010;
    wire [3:0] lut_438_select = {
                             in_data[120],
                             in_data[182],
                             in_data[334],
                             in_data[548]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b0001001100110011;
    wire [3:0] lut_439_select = {
                             in_data[199],
                             in_data[4],
                             in_data[18],
                             in_data[183]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b1000000011101101;
    wire [3:0] lut_440_select = {
                             in_data[158],
                             in_data[376],
                             in_data[116],
                             in_data[504]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b0000011100000111;
    wire [3:0] lut_441_select = {
                             in_data[415],
                             in_data[417],
                             in_data[527],
                             in_data[494]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b0011101100010000;
    wire [3:0] lut_442_select = {
                             in_data[530],
                             in_data[399],
                             in_data[352],
                             in_data[96]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1101010011110100;
    wire [3:0] lut_443_select = {
                             in_data[568],
                             in_data[275],
                             in_data[209],
                             in_data[127]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b1111001010110010;
    wire [3:0] lut_444_select = {
                             in_data[57],
                             in_data[86],
                             in_data[343],
                             in_data[406]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b0011111100101010;
    wire [3:0] lut_445_select = {
                             in_data[145],
                             in_data[64],
                             in_data[186],
                             in_data[22]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b0010111100001000;
    wire [3:0] lut_446_select = {
                             in_data[201],
                             in_data[160],
                             in_data[546],
                             in_data[413]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b0100010001011100;
    wire [3:0] lut_447_select = {
                             in_data[58],
                             in_data[383],
                             in_data[480],
                             in_data[342]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b1111100011100000;
    wire [3:0] lut_448_select = {
                             in_data[41],
                             in_data[78],
                             in_data[545],
                             in_data[374]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b0011111100110011;
    wire [3:0] lut_449_select = {
                             in_data[582],
                             in_data[172],
                             in_data[126],
                             in_data[102]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b0100110111111111;
    wire [3:0] lut_450_select = {
                             in_data[99],
                             in_data[423],
                             in_data[32],
                             in_data[164]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b0011101100101011;
    wire [3:0] lut_451_select = {
                             in_data[364],
                             in_data[139],
                             in_data[262],
                             in_data[265]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b1111011100010000;
    wire [3:0] lut_452_select = {
                             in_data[613],
                             in_data[1],
                             in_data[155],
                             in_data[299]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b1101110111011100;
    wire [3:0] lut_453_select = {
                             in_data[173],
                             in_data[10],
                             in_data[499],
                             in_data[69]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0010000010110011;
    wire [3:0] lut_454_select = {
                             in_data[431],
                             in_data[609],
                             in_data[384],
                             in_data[458]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b1100100011001100;
    wire [3:0] lut_455_select = {
                             in_data[106],
                             in_data[48],
                             in_data[216],
                             in_data[441]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b1101110111001100;
    wire [3:0] lut_456_select = {
                             in_data[240],
                             in_data[378],
                             in_data[427],
                             in_data[623]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b0111001101110111;
    wire [3:0] lut_457_select = {
                             in_data[101],
                             in_data[314],
                             in_data[303],
                             in_data[435]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b0010000010110000;
    wire [3:0] lut_458_select = {
                             in_data[393],
                             in_data[266],
                             in_data[189],
                             in_data[351]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b1111111100000000;
    wire [3:0] lut_459_select = {
                             in_data[462],
                             in_data[228],
                             in_data[570],
                             in_data[63]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b0101010101010111;
    wire [3:0] lut_460_select = {
                             in_data[614],
                             in_data[27],
                             in_data[354],
                             in_data[243]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b1101010111010101;
    wire [3:0] lut_461_select = {
                             in_data[624],
                             in_data[525],
                             in_data[484],
                             in_data[89]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b1110111011100000;
    wire [3:0] lut_462_select = {
                             in_data[481],
                             in_data[389],
                             in_data[146],
                             in_data[195]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b1111000011110100;
    wire [3:0] lut_463_select = {
                             in_data[516],
                             in_data[42],
                             in_data[198],
                             in_data[210]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b1000110000000000;
    wire [3:0] lut_464_select = {
                             in_data[402],
                             in_data[267],
                             in_data[236],
                             in_data[380]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b0010001010101010;
    wire [3:0] lut_465_select = {
                             in_data[282],
                             in_data[483],
                             in_data[79],
                             in_data[363]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b0000110101011111;
    wire [3:0] lut_466_select = {
                             in_data[249],
                             in_data[597],
                             in_data[340],
                             in_data[454]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1100110011001111;
    wire [3:0] lut_467_select = {
                             in_data[608],
                             in_data[226],
                             in_data[277],
                             in_data[241]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b0010101100111111;
    wire [3:0] lut_468_select = {
                             in_data[100],
                             in_data[124],
                             in_data[400],
                             in_data[50]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b0011000101110011;
    wire [3:0] lut_469_select = {
                             in_data[469],
                             in_data[17],
                             in_data[513],
                             in_data[118]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b0000111100001011;
    wire [3:0] lut_470_select = {
                             in_data[630],
                             in_data[111],
                             in_data[66],
                             in_data[75]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b0111001100110011;
    wire [3:0] lut_471_select = {
                             in_data[587],
                             in_data[439],
                             in_data[26],
                             in_data[391]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b0000111100001111;
    wire [3:0] lut_472_select = {
                             in_data[239],
                             in_data[612],
                             in_data[3],
                             in_data[167]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b1111111101010111;
    wire [3:0] lut_473_select = {
                             in_data[61],
                             in_data[412],
                             in_data[330],
                             in_data[252]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b0111011101110101;
    wire [3:0] lut_474_select = {
                             in_data[563],
                             in_data[531],
                             in_data[586],
                             in_data[325]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b1000100011101110;
    wire [3:0] lut_475_select = {
                             in_data[246],
                             in_data[135],
                             in_data[472],
                             in_data[33]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b0000111000001111;
    wire [3:0] lut_476_select = {
                             in_data[221],
                             in_data[87],
                             in_data[371],
                             in_data[577]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b1100110111011101;
    wire [3:0] lut_477_select = {
                             in_data[510],
                             in_data[457],
                             in_data[598],
                             in_data[593]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b1111000010000100;
    wire [3:0] lut_478_select = {
                             in_data[592],
                             in_data[373],
                             in_data[551],
                             in_data[543]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b0100010011111111;
    wire [3:0] lut_479_select = {
                             in_data[532],
                             in_data[72],
                             in_data[269],
                             in_data[178]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b0000010110111111;
    wire [3:0] lut_480_select = {
                             in_data[103],
                             in_data[294],
                             in_data[634],
                             in_data[472]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b1000000011101100;
    wire [3:0] lut_481_select = {
                             in_data[68],
                             in_data[444],
                             in_data[513],
                             in_data[332]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b0000100011001111;
    wire [3:0] lut_482_select = {
                             in_data[461],
                             in_data[46],
                             in_data[35],
                             in_data[88]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b1111000011111000;
    wire [3:0] lut_483_select = {
                             in_data[143],
                             in_data[504],
                             in_data[375],
                             in_data[39]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b0000111100001111;
    wire [3:0] lut_484_select = {
                             in_data[267],
                             in_data[601],
                             in_data[628],
                             in_data[414]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b1111001111110010;
    wire [3:0] lut_485_select = {
                             in_data[142],
                             in_data[200],
                             in_data[521],
                             in_data[223]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b0100111000000100;
    wire [3:0] lut_486_select = {
                             in_data[542],
                             in_data[44],
                             in_data[333],
                             in_data[576]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b0010001100100011;
    wire [3:0] lut_487_select = {
                             in_data[41],
                             in_data[522],
                             in_data[290],
                             in_data[323]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1111000101110000;
    wire [3:0] lut_488_select = {
                             in_data[297],
                             in_data[2],
                             in_data[562],
                             in_data[626]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b0111111100110111;
    wire [3:0] lut_489_select = {
                             in_data[558],
                             in_data[228],
                             in_data[439],
                             in_data[572]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b0001010100010111;
    wire [3:0] lut_490_select = {
                             in_data[420],
                             in_data[28],
                             in_data[604],
                             in_data[78]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b0000001001110011;
    wire [3:0] lut_491_select = {
                             in_data[496],
                             in_data[274],
                             in_data[411],
                             in_data[520]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b0010000000110011;
    wire [3:0] lut_492_select = {
                             in_data[292],
                             in_data[112],
                             in_data[340],
                             in_data[557]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b0000110011001111;
    wire [3:0] lut_493_select = {
                             in_data[239],
                             in_data[402],
                             in_data[624],
                             in_data[61]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b0001001100000001;
    wire [3:0] lut_494_select = {
                             in_data[413],
                             in_data[567],
                             in_data[91],
                             in_data[426]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b0000000011111111;
    wire [3:0] lut_495_select = {
                             in_data[531],
                             in_data[174],
                             in_data[328],
                             in_data[638]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b1011111110000010;
    wire [3:0] lut_496_select = {
                             in_data[145],
                             in_data[101],
                             in_data[373],
                             in_data[410]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b1101010011000100;
    wire [3:0] lut_497_select = {
                             in_data[178],
                             in_data[617],
                             in_data[519],
                             in_data[453]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b0111111101010111;
    wire [3:0] lut_498_select = {
                             in_data[72],
                             in_data[552],
                             in_data[443],
                             in_data[246]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b0000100011001110;
    wire [3:0] lut_499_select = {
                             in_data[425],
                             in_data[462],
                             in_data[157],
                             in_data[586]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b0000000000100010;
    wire [3:0] lut_500_select = {
                             in_data[129],
                             in_data[465],
                             in_data[484],
                             in_data[170]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b0001111100000001;
    wire [3:0] lut_501_select = {
                             in_data[321],
                             in_data[59],
                             in_data[302],
                             in_data[264]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b0000001100000111;
    wire [3:0] lut_502_select = {
                             in_data[283],
                             in_data[349],
                             in_data[573],
                             in_data[564]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b0010000110111011;
    wire [3:0] lut_503_select = {
                             in_data[151],
                             in_data[6],
                             in_data[155],
                             in_data[140]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b1101010011011101;
    wire [3:0] lut_504_select = {
                             in_data[296],
                             in_data[540],
                             in_data[547],
                             in_data[251]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b0010000011111111;
    wire [3:0] lut_505_select = {
                             in_data[190],
                             in_data[185],
                             in_data[368],
                             in_data[516]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b1011100011111010;
    wire [3:0] lut_506_select = {
                             in_data[153],
                             in_data[478],
                             in_data[172],
                             in_data[199]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b0011011100000000;
    wire [3:0] lut_507_select = {
                             in_data[236],
                             in_data[389],
                             in_data[249],
                             in_data[227]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b1111110011100000;
    wire [3:0] lut_508_select = {
                             in_data[127],
                             in_data[130],
                             in_data[337],
                             in_data[10]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b0000000011010101;
    wire [3:0] lut_509_select = {
                             in_data[204],
                             in_data[416],
                             in_data[448],
                             in_data[639]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b0101111100000101;
    wire [3:0] lut_510_select = {
                             in_data[355],
                             in_data[511],
                             in_data[554],
                             in_data[445]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0010000000110010;
    wire [3:0] lut_511_select = {
                             in_data[360],
                             in_data[109],
                             in_data[419],
                             in_data[0]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [15:0] lut_512_table = 16'b0001000100010001;
    wire [3:0] lut_512_select = {
                             in_data[73],
                             in_data[134],
                             in_data[481],
                             in_data[235]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [15:0] lut_513_table = 16'b1010000110000000;
    wire [3:0] lut_513_select = {
                             in_data[180],
                             in_data[238],
                             in_data[596],
                             in_data[5]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [15:0] lut_514_table = 16'b0100010001001111;
    wire [3:0] lut_514_select = {
                             in_data[629],
                             in_data[125],
                             in_data[428],
                             in_data[591]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [15:0] lut_515_table = 16'b0011000100110011;
    wire [3:0] lut_515_select = {
                             in_data[133],
                             in_data[118],
                             in_data[14],
                             in_data[255]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [15:0] lut_516_table = 16'b0101010100010000;
    wire [3:0] lut_516_select = {
                             in_data[363],
                             in_data[148],
                             in_data[300],
                             in_data[268]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [15:0] lut_517_table = 16'b1011101000001010;
    wire [3:0] lut_517_select = {
                             in_data[79],
                             in_data[231],
                             in_data[135],
                             in_data[21]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [15:0] lut_518_table = 16'b1111010011110101;
    wire [3:0] lut_518_select = {
                             in_data[146],
                             in_data[393],
                             in_data[34],
                             in_data[598]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [15:0] lut_519_table = 16'b1011101100101010;
    wire [3:0] lut_519_select = {
                             in_data[285],
                             in_data[19],
                             in_data[126],
                             in_data[526]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [15:0] lut_520_table = 16'b1111001100100000;
    wire [3:0] lut_520_select = {
                             in_data[560],
                             in_data[380],
                             in_data[354],
                             in_data[271]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [15:0] lut_521_table = 16'b1111111100001100;
    wire [3:0] lut_521_select = {
                             in_data[24],
                             in_data[430],
                             in_data[256],
                             in_data[501]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [15:0] lut_522_table = 16'b0011000100101010;
    wire [3:0] lut_522_select = {
                             in_data[429],
                             in_data[269],
                             in_data[571],
                             in_data[350]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [15:0] lut_523_table = 16'b1111111110000000;
    wire [3:0] lut_523_select = {
                             in_data[38],
                             in_data[523],
                             in_data[395],
                             in_data[463]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [15:0] lut_524_table = 16'b0001001100010101;
    wire [3:0] lut_524_select = {
                             in_data[440],
                             in_data[503],
                             in_data[74],
                             in_data[374]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [15:0] lut_525_table = 16'b0010001011111111;
    wire [3:0] lut_525_select = {
                             in_data[116],
                             in_data[376],
                             in_data[171],
                             in_data[635]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [15:0] lut_526_table = 16'b0101000001010000;
    wire [3:0] lut_526_select = {
                             in_data[92],
                             in_data[422],
                             in_data[114],
                             in_data[508]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [15:0] lut_527_table = 16'b1100111100000000;
    wire [3:0] lut_527_select = {
                             in_data[309],
                             in_data[3],
                             in_data[575],
                             in_data[442]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [15:0] lut_528_table = 16'b1010100010000000;
    wire [3:0] lut_528_select = {
                             in_data[110],
                             in_data[32],
                             in_data[154],
                             in_data[485]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [15:0] lut_529_table = 16'b1101110101000101;
    wire [3:0] lut_529_select = {
                             in_data[209],
                             in_data[330],
                             in_data[570],
                             in_data[213]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [15:0] lut_530_table = 16'b0100010011001111;
    wire [3:0] lut_530_select = {
                             in_data[315],
                             in_data[50],
                             in_data[275],
                             in_data[202]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [15:0] lut_531_table = 16'b1111001100110001;
    wire [3:0] lut_531_select = {
                             in_data[286],
                             in_data[122],
                             in_data[546],
                             in_data[351]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [15:0] lut_532_table = 16'b1111111101110011;
    wire [3:0] lut_532_select = {
                             in_data[131],
                             in_data[618],
                             in_data[208],
                             in_data[456]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [15:0] lut_533_table = 16'b0011010101110011;
    wire [3:0] lut_533_select = {
                             in_data[1],
                             in_data[466],
                             in_data[334],
                             in_data[359]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [15:0] lut_534_table = 16'b1011001011110000;
    wire [3:0] lut_534_select = {
                             in_data[207],
                             in_data[555],
                             in_data[600],
                             in_data[89]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [15:0] lut_535_table = 16'b1110110011101100;
    wire [3:0] lut_535_select = {
                             in_data[113],
                             in_data[587],
                             in_data[288],
                             in_data[121]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [15:0] lut_536_table = 16'b0101111101010000;
    wire [3:0] lut_536_select = {
                             in_data[270],
                             in_data[212],
                             in_data[347],
                             in_data[589]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [15:0] lut_537_table = 16'b1101000000000000;
    wire [3:0] lut_537_select = {
                             in_data[64],
                             in_data[424],
                             in_data[98],
                             in_data[167]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [15:0] lut_538_table = 16'b0111011100110010;
    wire [3:0] lut_538_select = {
                             in_data[336],
                             in_data[595],
                             in_data[406],
                             in_data[460]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [15:0] lut_539_table = 16'b0101110011001101;
    wire [3:0] lut_539_select = {
                             in_data[250],
                             in_data[631],
                             in_data[187],
                             in_data[450]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [15:0] lut_540_table = 16'b0000111100011111;
    wire [3:0] lut_540_select = {
                             in_data[47],
                             in_data[369],
                             in_data[509],
                             in_data[280]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [15:0] lut_541_table = 16'b0011000000110000;
    wire [3:0] lut_541_select = {
                             in_data[105],
                             in_data[473],
                             in_data[37],
                             in_data[175]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [15:0] lut_542_table = 16'b0101010011010101;
    wire [3:0] lut_542_select = {
                             in_data[408],
                             in_data[12],
                             in_data[353],
                             in_data[259]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [15:0] lut_543_table = 16'b0011001101111111;
    wire [3:0] lut_543_select = {
                             in_data[62],
                             in_data[470],
                             in_data[379],
                             in_data[124]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [15:0] lut_544_table = 16'b0000001000001111;
    wire [3:0] lut_544_select = {
                             in_data[561],
                             in_data[31],
                             in_data[317],
                             in_data[579]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [15:0] lut_545_table = 16'b0000010011001111;
    wire [3:0] lut_545_select = {
                             in_data[335],
                             in_data[273],
                             in_data[99],
                             in_data[211]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [15:0] lut_546_table = 16'b0111111100001100;
    wire [3:0] lut_546_select = {
                             in_data[582],
                             in_data[348],
                             in_data[100],
                             in_data[468]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [15:0] lut_547_table = 16'b0011000110111111;
    wire [3:0] lut_547_select = {
                             in_data[489],
                             in_data[569],
                             in_data[137],
                             in_data[198]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [15:0] lut_548_table = 16'b0011001100110011;
    wire [3:0] lut_548_select = {
                             in_data[253],
                             in_data[104],
                             in_data[342],
                             in_data[486]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [15:0] lut_549_table = 16'b0011000000110000;
    wire [3:0] lut_549_select = {
                             in_data[475],
                             in_data[293],
                             in_data[82],
                             in_data[610]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [15:0] lut_550_table = 16'b0101010001000100;
    wire [3:0] lut_550_select = {
                             in_data[195],
                             in_data[188],
                             in_data[563],
                             in_data[417]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [15:0] lut_551_table = 16'b0000111011001111;
    wire [3:0] lut_551_select = {
                             in_data[344],
                             in_data[479],
                             in_data[447],
                             in_data[320]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [15:0] lut_552_table = 16'b0000101100111011;
    wire [3:0] lut_552_select = {
                             in_data[243],
                             in_data[95],
                             in_data[318],
                             in_data[97]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [15:0] lut_553_table = 16'b0100010111111111;
    wire [3:0] lut_553_select = {
                             in_data[26],
                             in_data[13],
                             in_data[177],
                             in_data[107]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [15:0] lut_554_table = 16'b1100111011001111;
    wire [3:0] lut_554_select = {
                             in_data[36],
                             in_data[83],
                             in_data[229],
                             in_data[42]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [15:0] lut_555_table = 16'b0001010001010101;
    wire [3:0] lut_555_select = {
                             in_data[240],
                             in_data[559],
                             in_data[291],
                             in_data[597]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [15:0] lut_556_table = 16'b1000111010101111;
    wire [3:0] lut_556_select = {
                             in_data[40],
                             in_data[396],
                             in_data[609],
                             in_data[619]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [15:0] lut_557_table = 16'b0000100000001100;
    wire [3:0] lut_557_select = {
                             in_data[196],
                             in_data[605],
                             in_data[625],
                             in_data[482]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [15:0] lut_558_table = 16'b1011101100100010;
    wire [3:0] lut_558_select = {
                             in_data[515],
                             in_data[96],
                             in_data[169],
                             in_data[537]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [15:0] lut_559_table = 16'b0000110100000100;
    wire [3:0] lut_559_select = {
                             in_data[272],
                             in_data[7],
                             in_data[316],
                             in_data[592]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [15:0] lut_560_table = 16'b0000110000001101;
    wire [3:0] lut_560_select = {
                             in_data[329],
                             in_data[299],
                             in_data[49],
                             in_data[459]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [15:0] lut_561_table = 16'b0101111101011111;
    wire [3:0] lut_561_select = {
                             in_data[434],
                             in_data[54],
                             in_data[277],
                             in_data[517]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [15:0] lut_562_table = 16'b1111111111101000;
    wire [3:0] lut_562_select = {
                             in_data[580],
                             in_data[584],
                             in_data[65],
                             in_data[52]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [15:0] lut_563_table = 16'b1111111100111111;
    wire [3:0] lut_563_select = {
                             in_data[630],
                             in_data[585],
                             in_data[616],
                             in_data[77]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [15:0] lut_564_table = 16'b1111111110001000;
    wire [3:0] lut_564_select = {
                             in_data[67],
                             in_data[487],
                             in_data[18],
                             in_data[115]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [15:0] lut_565_table = 16'b1000111011001111;
    wire [3:0] lut_565_select = {
                             in_data[132],
                             in_data[70],
                             in_data[76],
                             in_data[588]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [15:0] lut_566_table = 16'b0010000011111010;
    wire [3:0] lut_566_select = {
                             in_data[224],
                             in_data[464],
                             in_data[282],
                             in_data[310]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [15:0] lut_567_table = 16'b0101000001000100;
    wire [3:0] lut_567_select = {
                             in_data[533],
                             in_data[136],
                             in_data[544],
                             in_data[254]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [15:0] lut_568_table = 16'b1010000010101000;
    wire [3:0] lut_568_select = {
                             in_data[409],
                             in_data[191],
                             in_data[203],
                             in_data[599]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [15:0] lut_569_table = 16'b0101111100000101;
    wire [3:0] lut_569_select = {
                             in_data[502],
                             in_data[433],
                             in_data[232],
                             in_data[25]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [15:0] lut_570_table = 16'b0101111101011111;
    wire [3:0] lut_570_select = {
                             in_data[357],
                             in_data[623],
                             in_data[390],
                             in_data[632]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [15:0] lut_571_table = 16'b0100010001010100;
    wire [3:0] lut_571_select = {
                             in_data[308],
                             in_data[452],
                             in_data[493],
                             in_data[483]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [15:0] lut_572_table = 16'b0000101010101011;
    wire [3:0] lut_572_select = {
                             in_data[614],
                             in_data[367],
                             in_data[119],
                             in_data[471]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [15:0] lut_573_table = 16'b0011001000100010;
    wire [3:0] lut_573_select = {
                             in_data[162],
                             in_data[613],
                             in_data[222],
                             in_data[248]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [15:0] lut_574_table = 16'b0001001101011111;
    wire [3:0] lut_574_select = {
                             in_data[276],
                             in_data[602],
                             in_data[166],
                             in_data[405]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [15:0] lut_575_table = 16'b1011001111110011;
    wire [3:0] lut_575_select = {
                             in_data[438],
                             in_data[45],
                             in_data[548],
                             in_data[492]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [15:0] lut_576_table = 16'b1111111100000111;
    wire [3:0] lut_576_select = {
                             in_data[633],
                             in_data[365],
                             in_data[193],
                             in_data[149]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [15:0] lut_577_table = 16'b1111101100100011;
    wire [3:0] lut_577_select = {
                             in_data[362],
                             in_data[120],
                             in_data[358],
                             in_data[205]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [15:0] lut_578_table = 16'b0101011101010111;
    wire [3:0] lut_578_select = {
                             in_data[9],
                             in_data[556],
                             in_data[201],
                             in_data[301]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [15:0] lut_579_table = 16'b1010111010101010;
    wire [3:0] lut_579_select = {
                             in_data[566],
                             in_data[455],
                             in_data[234],
                             in_data[152]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [15:0] lut_580_table = 16'b1110111011001010;
    wire [3:0] lut_580_select = {
                             in_data[314],
                             in_data[261],
                             in_data[22],
                             in_data[361]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [15:0] lut_581_table = 16'b0001001111111111;
    wire [3:0] lut_581_select = {
                             in_data[30],
                             in_data[27],
                             in_data[467],
                             in_data[128]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [15:0] lut_582_table = 16'b0011101100101011;
    wire [3:0] lut_582_select = {
                             in_data[245],
                             in_data[55],
                             in_data[304],
                             in_data[63]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [15:0] lut_583_table = 16'b1010100010101000;
    wire [3:0] lut_583_select = {
                             in_data[33],
                             in_data[477],
                             in_data[322],
                             in_data[525]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [15:0] lut_584_table = 16'b1100111100001000;
    wire [3:0] lut_584_select = {
                             in_data[303],
                             in_data[512],
                             in_data[217],
                             in_data[106]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [15:0] lut_585_table = 16'b0000111100001010;
    wire [3:0] lut_585_select = {
                             in_data[266],
                             in_data[494],
                             in_data[221],
                             in_data[530]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [15:0] lut_586_table = 16'b0000111100001111;
    wire [3:0] lut_586_select = {
                             in_data[325],
                             in_data[446],
                             in_data[506],
                             in_data[53]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [15:0] lut_587_table = 16'b1100110011001111;
    wire [3:0] lut_587_select = {
                             in_data[392],
                             in_data[23],
                             in_data[451],
                             in_data[58]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [15:0] lut_588_table = 16'b1010111100001011;
    wire [3:0] lut_588_select = {
                             in_data[535],
                             in_data[305],
                             in_data[192],
                             in_data[138]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [15:0] lut_589_table = 16'b1111111100000101;
    wire [3:0] lut_589_select = {
                             in_data[182],
                             in_data[608],
                             in_data[534],
                             in_data[427]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [15:0] lut_590_table = 16'b0000000001110111;
    wire [3:0] lut_590_select = {
                             in_data[225],
                             in_data[284],
                             in_data[394],
                             in_data[524]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [15:0] lut_591_table = 16'b1111001111110000;
    wire [3:0] lut_591_select = {
                             in_data[326],
                             in_data[345],
                             in_data[421],
                             in_data[289]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [15:0] lut_592_table = 16'b1111001011110010;
    wire [3:0] lut_592_select = {
                             in_data[536],
                             in_data[144],
                             in_data[60],
                             in_data[622]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [15:0] lut_593_table = 16'b1111010101010000;
    wire [3:0] lut_593_select = {
                             in_data[539],
                             in_data[183],
                             in_data[435],
                             in_data[577]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [15:0] lut_594_table = 16'b0000010101111111;
    wire [3:0] lut_594_select = {
                             in_data[84],
                             in_data[403],
                             in_data[313],
                             in_data[385]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [15:0] lut_595_table = 16'b1111011101110000;
    wire [3:0] lut_595_select = {
                             in_data[527],
                             in_data[415],
                             in_data[543],
                             in_data[499]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [15:0] lut_596_table = 16'b1111010001100000;
    wire [3:0] lut_596_select = {
                             in_data[397],
                             in_data[75],
                             in_data[287],
                             in_data[71]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [15:0] lut_597_table = 16'b0000010111011111;
    wire [3:0] lut_597_select = {
                             in_data[510],
                             in_data[457],
                             in_data[189],
                             in_data[168]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [15:0] lut_598_table = 16'b0000010111010101;
    wire [3:0] lut_598_select = {
                             in_data[158],
                             in_data[352],
                             in_data[449],
                             in_data[164]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [15:0] lut_599_table = 16'b0100010011000100;
    wire [3:0] lut_599_select = {
                             in_data[431],
                             in_data[165],
                             in_data[549],
                             in_data[176]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [15:0] lut_600_table = 16'b1000111000001100;
    wire [3:0] lut_600_select = {
                             in_data[279],
                             in_data[495],
                             in_data[377],
                             in_data[491]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [15:0] lut_601_table = 16'b1000100011111011;
    wire [3:0] lut_601_select = {
                             in_data[8],
                             in_data[87],
                             in_data[480],
                             in_data[338]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [15:0] lut_602_table = 16'b0011000100110001;
    wire [3:0] lut_602_select = {
                             in_data[505],
                             in_data[565],
                             in_data[391],
                             in_data[43]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [15:0] lut_603_table = 16'b1110111011101010;
    wire [3:0] lut_603_select = {
                             in_data[545],
                             in_data[156],
                             in_data[159],
                             in_data[603]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [15:0] lut_604_table = 16'b0101010001010101;
    wire [3:0] lut_604_select = {
                             in_data[214],
                             in_data[20],
                             in_data[139],
                             in_data[219]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [15:0] lut_605_table = 16'b1010000011110000;
    wire [3:0] lut_605_select = {
                             in_data[111],
                             in_data[161],
                             in_data[606],
                             in_data[11]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [15:0] lut_606_table = 16'b1010001011111111;
    wire [3:0] lut_606_select = {
                             in_data[102],
                             in_data[295],
                             in_data[568],
                             in_data[615]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [15:0] lut_607_table = 16'b0010000100110001;
    wire [3:0] lut_607_select = {
                             in_data[147],
                             in_data[381],
                             in_data[339],
                             in_data[436]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [15:0] lut_608_table = 16'b1010101011111111;
    wire [3:0] lut_608_select = {
                             in_data[230],
                             in_data[260],
                             in_data[108],
                             in_data[94]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [15:0] lut_609_table = 16'b1111011111010000;
    wire [3:0] lut_609_select = {
                             in_data[611],
                             in_data[233],
                             in_data[593],
                             in_data[364]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [15:0] lut_610_table = 16'b1111110100000000;
    wire [3:0] lut_610_select = {
                             in_data[578],
                             in_data[197],
                             in_data[312],
                             in_data[514]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [15:0] lut_611_table = 16'b0010101000101010;
    wire [3:0] lut_611_select = {
                             in_data[319],
                             in_data[226],
                             in_data[636],
                             in_data[244]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [15:0] lut_612_table = 16'b1011001010101000;
    wire [3:0] lut_612_select = {
                             in_data[574],
                             in_data[29],
                             in_data[306],
                             in_data[551]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [15:0] lut_613_table = 16'b0000000010001110;
    wire [3:0] lut_613_select = {
                             in_data[437],
                             in_data[404],
                             in_data[343],
                             in_data[86]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [15:0] lut_614_table = 16'b1000101010011011;
    wire [3:0] lut_614_select = {
                             in_data[454],
                             in_data[194],
                             in_data[160],
                             in_data[507]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [15:0] lut_615_table = 16'b0011111100011111;
    wire [3:0] lut_615_select = {
                             in_data[553],
                             in_data[81],
                             in_data[93],
                             in_data[423]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [15:0] lut_616_table = 16'b0101111100000000;
    wire [3:0] lut_616_select = {
                             in_data[418],
                             in_data[383],
                             in_data[583],
                             in_data[141]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [15:0] lut_617_table = 16'b1011101110001011;
    wire [3:0] lut_617_select = {
                             in_data[298],
                             in_data[15],
                             in_data[621],
                             in_data[220]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [15:0] lut_618_table = 16'b0000101000101111;
    wire [3:0] lut_618_select = {
                             in_data[637],
                             in_data[66],
                             in_data[432],
                             in_data[627]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [15:0] lut_619_table = 16'b0000000011010101;
    wire [3:0] lut_619_select = {
                             in_data[179],
                             in_data[206],
                             in_data[371],
                             in_data[163]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [15:0] lut_620_table = 16'b1100111111001111;
    wire [3:0] lut_620_select = {
                             in_data[378],
                             in_data[529],
                             in_data[400],
                             in_data[497]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [15:0] lut_621_table = 16'b1101010011110100;
    wire [3:0] lut_621_select = {
                             in_data[458],
                             in_data[384],
                             in_data[370],
                             in_data[184]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [15:0] lut_622_table = 16'b1011101011111011;
    wire [3:0] lut_622_select = {
                             in_data[210],
                             in_data[56],
                             in_data[69],
                             in_data[518]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [15:0] lut_623_table = 16'b1010001100101011;
    wire [3:0] lut_623_select = {
                             in_data[469],
                             in_data[150],
                             in_data[117],
                             in_data[247]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [15:0] lut_624_table = 16'b0001001101010101;
    wire [3:0] lut_624_select = {
                             in_data[538],
                             in_data[181],
                             in_data[16],
                             in_data[281]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [15:0] lut_625_table = 16'b1111110001000000;
    wire [3:0] lut_625_select = {
                             in_data[257],
                             in_data[242],
                             in_data[237],
                             in_data[216]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [15:0] lut_626_table = 16'b0011111100001111;
    wire [3:0] lut_626_select = {
                             in_data[265],
                             in_data[341],
                             in_data[17],
                             in_data[366]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [15:0] lut_627_table = 16'b0101110101011111;
    wire [3:0] lut_627_select = {
                             in_data[476],
                             in_data[241],
                             in_data[48],
                             in_data[331]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [15:0] lut_628_table = 16'b0100010011001101;
    wire [3:0] lut_628_select = {
                             in_data[51],
                             in_data[356],
                             in_data[57],
                             in_data[324]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [15:0] lut_629_table = 16'b0000000100111111;
    wire [3:0] lut_629_select = {
                             in_data[401],
                             in_data[528],
                             in_data[620],
                             in_data[412]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [15:0] lut_630_table = 16'b0010001000001010;
    wire [3:0] lut_630_select = {
                             in_data[488],
                             in_data[4],
                             in_data[541],
                             in_data[590]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [15:0] lut_631_table = 16'b0011001010110010;
    wire [3:0] lut_631_select = {
                             in_data[581],
                             in_data[80],
                             in_data[388],
                             in_data[386]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [15:0] lut_632_table = 16'b1111000011000000;
    wire [3:0] lut_632_select = {
                             in_data[123],
                             in_data[173],
                             in_data[594],
                             in_data[490]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [15:0] lut_633_table = 16'b1000100011101010;
    wire [3:0] lut_633_select = {
                             in_data[252],
                             in_data[498],
                             in_data[307],
                             in_data[215]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [15:0] lut_634_table = 16'b0010101000100011;
    wire [3:0] lut_634_select = {
                             in_data[607],
                             in_data[186],
                             in_data[327],
                             in_data[372]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [15:0] lut_635_table = 16'b0111111100000101;
    wire [3:0] lut_635_select = {
                             in_data[398],
                             in_data[311],
                             in_data[612],
                             in_data[441]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [15:0] lut_636_table = 16'b0100010101000101;
    wire [3:0] lut_636_select = {
                             in_data[278],
                             in_data[85],
                             in_data[382],
                             in_data[474]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [15:0] lut_637_table = 16'b0101111100000101;
    wire [3:0] lut_637_select = {
                             in_data[263],
                             in_data[500],
                             in_data[218],
                             in_data[532]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [15:0] lut_638_table = 16'b0000011100000000;
    wire [3:0] lut_638_select = {
                             in_data[550],
                             in_data[407],
                             in_data[387],
                             in_data[90]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [15:0] lut_639_table = 16'b0000100000111111;
    wire [3:0] lut_639_select = {
                             in_data[258],
                             in_data[399],
                             in_data[346],
                             in_data[262]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub4
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        639:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        639:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub4_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub4_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub4_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [639:0]  in_data,
            output wire [639:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1101000011111100;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b0000000001010111;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b0000101110111111;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1111000011111111;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b1111110101010000;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1111010100110000;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b1011001011111011;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b0111000100010000;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b0101110111010101;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b0101111101011110;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b1010111100001011;
    wire [3:0] lut_10_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b1111111111010000;
    wire [3:0] lut_11_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b0111001011110010;
    wire [3:0] lut_12_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0000001100111111;
    wire [3:0] lut_13_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0111000111110011;
    wire [3:0] lut_14_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b0000011100111111;
    wire [3:0] lut_15_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b0000110000111111;
    wire [3:0] lut_16_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b1100110011000100;
    wire [3:0] lut_17_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0010001100111011;
    wire [3:0] lut_18_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b0000000010111011;
    wire [3:0] lut_19_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0000000011101111;
    wire [3:0] lut_20_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b0001011100000101;
    wire [3:0] lut_21_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b1111011111110001;
    wire [3:0] lut_22_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0000110011001110;
    wire [3:0] lut_23_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1111111111110100;
    wire [3:0] lut_24_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0011000000010000;
    wire [3:0] lut_25_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b0101111101010101;
    wire [3:0] lut_26_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1111111100110000;
    wire [3:0] lut_27_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b0011001100000000;
    wire [3:0] lut_28_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b0000010100010111;
    wire [3:0] lut_29_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b0000010001010101;
    wire [3:0] lut_30_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1011111111101110;
    wire [3:0] lut_31_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1011001100110010;
    wire [3:0] lut_32_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b1111010101000000;
    wire [3:0] lut_33_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1111011111110001;
    wire [3:0] lut_34_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1000101010101010;
    wire [3:0] lut_35_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b0000000011001000;
    wire [3:0] lut_36_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b1110111010001110;
    wire [3:0] lut_37_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b0100010001000100;
    wire [3:0] lut_38_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0101010011011101;
    wire [3:0] lut_39_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b0111111101010101;
    wire [3:0] lut_40_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b0000000000000011;
    wire [3:0] lut_41_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b0010101000000000;
    wire [3:0] lut_42_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0011001100110011;
    wire [3:0] lut_43_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b0000010100010111;
    wire [3:0] lut_44_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b1010100000000000;
    wire [3:0] lut_45_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b1101000011010000;
    wire [3:0] lut_46_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b1101010001000000;
    wire [3:0] lut_47_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b0011001011110011;
    wire [3:0] lut_48_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b0011001000110000;
    wire [3:0] lut_49_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b1111111111110001;
    wire [3:0] lut_50_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b0000111100001111;
    wire [3:0] lut_51_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1010111000000000;
    wire [3:0] lut_52_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b0111000100010000;
    wire [3:0] lut_53_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b1101110101010100;
    wire [3:0] lut_54_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b1010100010001000;
    wire [3:0] lut_55_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b0000010101011111;
    wire [3:0] lut_56_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b0000000010101010;
    wire [3:0] lut_57_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b0000110110001110;
    wire [3:0] lut_58_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b1011101010110010;
    wire [3:0] lut_59_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b0001000101010101;
    wire [3:0] lut_60_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b0001001100000111;
    wire [3:0] lut_61_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b0111000100000000;
    wire [3:0] lut_62_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b0000000101011111;
    wire [3:0] lut_63_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b0000111111111111;
    wire [3:0] lut_64_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b1110111000001110;
    wire [3:0] lut_65_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b0010000010110010;
    wire [3:0] lut_66_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b0100110100000000;
    wire [3:0] lut_67_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b0101010011011100;
    wire [3:0] lut_68_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b1110000011100000;
    wire [3:0] lut_69_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b0010001000100010;
    wire [3:0] lut_70_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0101000101110001;
    wire [3:0] lut_71_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b0000111010101111;
    wire [3:0] lut_72_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b0010111000101011;
    wire [3:0] lut_73_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0111010101010101;
    wire [3:0] lut_74_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b0111000101110101;
    wire [3:0] lut_75_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0100010101000101;
    wire [3:0] lut_76_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b1111001111110010;
    wire [3:0] lut_77_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b1111110111010100;
    wire [3:0] lut_78_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b0101000100000001;
    wire [3:0] lut_79_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b0011000001110001;
    wire [3:0] lut_80_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b1111110001010000;
    wire [3:0] lut_81_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1111111100001111;
    wire [3:0] lut_82_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b0000111010001111;
    wire [3:0] lut_83_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b0101111100000100;
    wire [3:0] lut_84_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b0000010101010111;
    wire [3:0] lut_85_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b1101010101000101;
    wire [3:0] lut_86_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b1011001011111011;
    wire [3:0] lut_87_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b0101000001110011;
    wire [3:0] lut_88_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b0001010101010101;
    wire [3:0] lut_89_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1000111100001011;
    wire [3:0] lut_90_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b1111000011111100;
    wire [3:0] lut_91_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1111110011111100;
    wire [3:0] lut_92_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0000110010001111;
    wire [3:0] lut_93_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b0000000100110011;
    wire [3:0] lut_94_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b0100010101000100;
    wire [3:0] lut_95_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1011101100100010;
    wire [3:0] lut_96_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b1111111101000101;
    wire [3:0] lut_97_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1111101000100010;
    wire [3:0] lut_98_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b0000101010101111;
    wire [3:0] lut_99_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1101110111011100;
    wire [3:0] lut_100_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b0011000011111111;
    wire [3:0] lut_101_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b0010001010111111;
    wire [3:0] lut_102_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1000100011101110;
    wire [3:0] lut_103_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b1110100000000000;
    wire [3:0] lut_104_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1011101010111011;
    wire [3:0] lut_105_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b1110100011111110;
    wire [3:0] lut_106_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b1111001000000000;
    wire [3:0] lut_107_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b0001111101111111;
    wire [3:0] lut_108_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b0000110011001100;
    wire [3:0] lut_109_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b0000001100111111;
    wire [3:0] lut_110_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000100000001110;
    wire [3:0] lut_111_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b1011101110110011;
    wire [3:0] lut_112_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b1100000011011100;
    wire [3:0] lut_113_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1111010011110101;
    wire [3:0] lut_114_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0101000011010100;
    wire [3:0] lut_115_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b1111111011101100;
    wire [3:0] lut_116_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b1111100011100000;
    wire [3:0] lut_117_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1101010011000000;
    wire [3:0] lut_118_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b1111111100100010;
    wire [3:0] lut_119_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b0000111010101111;
    wire [3:0] lut_120_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b1111111100000010;
    wire [3:0] lut_121_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b1011111100101111;
    wire [3:0] lut_122_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b0000110000001100;
    wire [3:0] lut_123_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b0000000001110011;
    wire [3:0] lut_124_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b1111111010101010;
    wire [3:0] lut_125_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b1111101100110011;
    wire [3:0] lut_126_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0000000010001010;
    wire [3:0] lut_127_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b1111001110110011;
    wire [3:0] lut_128_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b1010000011111011;
    wire [3:0] lut_129_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b1111101100100010;
    wire [3:0] lut_130_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b1111111111110001;
    wire [3:0] lut_131_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b1011111110101010;
    wire [3:0] lut_132_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0101111111010101;
    wire [3:0] lut_133_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b0111010100010000;
    wire [3:0] lut_134_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b0001000000110000;
    wire [3:0] lut_135_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b0000000100010111;
    wire [3:0] lut_136_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b1111110111110100;
    wire [3:0] lut_137_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b0111000101110001;
    wire [3:0] lut_138_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b1100111101001101;
    wire [3:0] lut_139_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b0000111111111111;
    wire [3:0] lut_140_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b0100010011011111;
    wire [3:0] lut_141_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b1011000010110010;
    wire [3:0] lut_142_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0010101000100010;
    wire [3:0] lut_143_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b0011000000110000;
    wire [3:0] lut_144_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1110111010000000;
    wire [3:0] lut_145_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b0011000010110000;
    wire [3:0] lut_146_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0010001101110111;
    wire [3:0] lut_147_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b0011001000110010;
    wire [3:0] lut_148_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b0011101110111011;
    wire [3:0] lut_149_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b0000010100001111;
    wire [3:0] lut_150_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b0100111111011111;
    wire [3:0] lut_151_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b1110111011001000;
    wire [3:0] lut_152_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1111110011010100;
    wire [3:0] lut_153_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0011011100100111;
    wire [3:0] lut_154_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b0000000010101000;
    wire [3:0] lut_155_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b0011000001110000;
    wire [3:0] lut_156_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b1110111110001000;
    wire [3:0] lut_157_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b0111000011110001;
    wire [3:0] lut_158_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b0010101100101111;
    wire [3:0] lut_159_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b0101000111110111;
    wire [3:0] lut_160_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b0001000100110011;
    wire [3:0] lut_161_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1101010101000000;
    wire [3:0] lut_162_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b0101111100000111;
    wire [3:0] lut_163_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b0000001000001011;
    wire [3:0] lut_164_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b1000100011101110;
    wire [3:0] lut_165_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b0000110100000000;
    wire [3:0] lut_166_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b0111011100010001;
    wire [3:0] lut_167_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b1101010111010100;
    wire [3:0] lut_168_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b1010100010001000;
    wire [3:0] lut_169_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b1101000011110100;
    wire [3:0] lut_170_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b1000000011111101;
    wire [3:0] lut_171_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b0001000101010101;
    wire [3:0] lut_172_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b0000011101111111;
    wire [3:0] lut_173_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b0011000001110010;
    wire [3:0] lut_174_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1000100010000000;
    wire [3:0] lut_175_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b1111001111010000;
    wire [3:0] lut_176_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b1000110010001110;
    wire [3:0] lut_177_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b0110111100100010;
    wire [3:0] lut_178_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b1110100011111110;
    wire [3:0] lut_179_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b1000100010001000;
    wire [3:0] lut_180_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b0001011100000001;
    wire [3:0] lut_181_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b1000100011001111;
    wire [3:0] lut_182_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b0000110001001111;
    wire [3:0] lut_183_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b0000000000001011;
    wire [3:0] lut_184_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b0111000100010000;
    wire [3:0] lut_185_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b0111101100010000;
    wire [3:0] lut_186_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b1101110111011101;
    wire [3:0] lut_187_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b0101110101011111;
    wire [3:0] lut_188_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b1011101100100011;
    wire [3:0] lut_189_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b1101010001000000;
    wire [3:0] lut_190_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b1110111000001100;
    wire [3:0] lut_191_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b1100110011001101;
    wire [3:0] lut_192_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b0000101011111111;
    wire [3:0] lut_193_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0000111000001101;
    wire [3:0] lut_194_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b1000111110001110;
    wire [3:0] lut_195_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b1100010011010100;
    wire [3:0] lut_196_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b1010111010101110;
    wire [3:0] lut_197_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b0110000011110010;
    wire [3:0] lut_198_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b1101110101011101;
    wire [3:0] lut_199_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b0000000011110010;
    wire [3:0] lut_200_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b1111010111010100;
    wire [3:0] lut_201_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b1010101000000000;
    wire [3:0] lut_202_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b0000101010101110;
    wire [3:0] lut_203_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b1111101010111000;
    wire [3:0] lut_204_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b0001011111111111;
    wire [3:0] lut_205_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b0111111100000011;
    wire [3:0] lut_206_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b0101010101000100;
    wire [3:0] lut_207_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1000111100000100;
    wire [3:0] lut_208_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b1100111101001110;
    wire [3:0] lut_209_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b0000111010001111;
    wire [3:0] lut_210_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b1011111100001111;
    wire [3:0] lut_211_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b0011001100110011;
    wire [3:0] lut_212_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b0000010001011101;
    wire [3:0] lut_213_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1111110111010100;
    wire [3:0] lut_214_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b1100100010100000;
    wire [3:0] lut_215_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b1010101010100000;
    wire [3:0] lut_216_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b0111111100000101;
    wire [3:0] lut_217_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b1111111100010000;
    wire [3:0] lut_218_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b0100010100000100;
    wire [3:0] lut_219_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b0001000001110011;
    wire [3:0] lut_220_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b0010001000101011;
    wire [3:0] lut_221_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b0111000100000000;
    wire [3:0] lut_222_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1110110011001100;
    wire [3:0] lut_223_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b1111000000000000;
    wire [3:0] lut_224_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b1100111100001110;
    wire [3:0] lut_225_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1011001010110010;
    wire [3:0] lut_226_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b1011000011110011;
    wire [3:0] lut_227_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b1111001100100010;
    wire [3:0] lut_228_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b1110101010000000;
    wire [3:0] lut_229_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b0000010011011101;
    wire [3:0] lut_230_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b0010111100010001;
    wire [3:0] lut_231_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b0100010011001100;
    wire [3:0] lut_232_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b1100000011101100;
    wire [3:0] lut_233_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b0000100010001110;
    wire [3:0] lut_234_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b0010101010101011;
    wire [3:0] lut_235_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b0101110111111111;
    wire [3:0] lut_236_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b0011000011110111;
    wire [3:0] lut_237_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b0000001010101010;
    wire [3:0] lut_238_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0000111100001110;
    wire [3:0] lut_239_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b0111000101110001;
    wire [3:0] lut_240_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b0000111110001111;
    wire [3:0] lut_241_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b0000111101000101;
    wire [3:0] lut_242_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b0000100010001000;
    wire [3:0] lut_243_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b1110000011111010;
    wire [3:0] lut_244_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b1110101011101000;
    wire [3:0] lut_245_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b0101111100001010;
    wire [3:0] lut_246_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b1100111100001100;
    wire [3:0] lut_247_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b0011001111110111;
    wire [3:0] lut_248_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b1111111011100000;
    wire [3:0] lut_249_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b0011000111110111;
    wire [3:0] lut_250_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b1110000011110100;
    wire [3:0] lut_251_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b0010101100001000;
    wire [3:0] lut_252_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b1000111010001111;
    wire [3:0] lut_253_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b1110111011101000;
    wire [3:0] lut_254_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b0001001100000001;
    wire [3:0] lut_255_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b1011101100110011;
    wire [3:0] lut_256_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b1101111101001101;
    wire [3:0] lut_257_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b0001011100110111;
    wire [3:0] lut_258_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b1100111011101111;
    wire [3:0] lut_259_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b1111000011110100;
    wire [3:0] lut_260_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b0010101010111011;
    wire [3:0] lut_261_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b1101110101000000;
    wire [3:0] lut_262_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b1110010011111110;
    wire [3:0] lut_263_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b0001001100111111;
    wire [3:0] lut_264_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b1100010011111101;
    wire [3:0] lut_265_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1111101011111010;
    wire [3:0] lut_266_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b0001011100010111;
    wire [3:0] lut_267_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1100010000000000;
    wire [3:0] lut_268_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0111011101110101;
    wire [3:0] lut_269_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b0000001100111111;
    wire [3:0] lut_270_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b0100010001001101;
    wire [3:0] lut_271_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b0100110101011111;
    wire [3:0] lut_272_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b0011111100000011;
    wire [3:0] lut_273_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b1111111100110011;
    wire [3:0] lut_274_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b1100110011000100;
    wire [3:0] lut_275_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b1111101011101110;
    wire [3:0] lut_276_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b1110110010001000;
    wire [3:0] lut_277_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b0010001010111111;
    wire [3:0] lut_278_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b0000010001010101;
    wire [3:0] lut_279_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b1100111111001111;
    wire [3:0] lut_280_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b1111101010101000;
    wire [3:0] lut_281_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b0100010011001101;
    wire [3:0] lut_282_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b1111000011111010;
    wire [3:0] lut_283_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b1100111111001100;
    wire [3:0] lut_284_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b0000110000001111;
    wire [3:0] lut_285_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b0000111000001110;
    wire [3:0] lut_286_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b0010000010101011;
    wire [3:0] lut_287_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b1111010101010000;
    wire [3:0] lut_288_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b0100110001011101;
    wire [3:0] lut_289_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b0010001100100010;
    wire [3:0] lut_290_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b0000100010001110;
    wire [3:0] lut_291_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b1011101110101011;
    wire [3:0] lut_292_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b0010000000100010;
    wire [3:0] lut_293_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1100111111001101;
    wire [3:0] lut_294_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b1101110011000100;
    wire [3:0] lut_295_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b1111100011111100;
    wire [3:0] lut_296_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b1111110111110101;
    wire [3:0] lut_297_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b1000111010001110;
    wire [3:0] lut_298_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b0010000010110000;
    wire [3:0] lut_299_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b0101000100010001;
    wire [3:0] lut_300_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b1111110011110100;
    wire [3:0] lut_301_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b1100111101001100;
    wire [3:0] lut_302_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b1010001100100000;
    wire [3:0] lut_303_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b1000111011001111;
    wire [3:0] lut_304_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b1000100010000000;
    wire [3:0] lut_305_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b1100111111001100;
    wire [3:0] lut_306_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b0010001101110111;
    wire [3:0] lut_307_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b0001010001111111;
    wire [3:0] lut_308_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b1101000011111000;
    wire [3:0] lut_309_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b0101011100000001;
    wire [3:0] lut_310_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b1111101010100000;
    wire [3:0] lut_311_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1111111010001000;
    wire [3:0] lut_312_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b1101110111010100;
    wire [3:0] lut_313_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b1100111110001000;
    wire [3:0] lut_314_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b1111000100110000;
    wire [3:0] lut_315_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b1000111010101111;
    wire [3:0] lut_316_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b0011000100110001;
    wire [3:0] lut_317_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0011000011110011;
    wire [3:0] lut_318_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b0000001100010111;
    wire [3:0] lut_319_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b0001000100110111;
    wire [3:0] lut_320_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0001000011110001;
    wire [3:0] lut_321_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b1000101010101111;
    wire [3:0] lut_322_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b1111111100000001;
    wire [3:0] lut_323_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b0000101000001111;
    wire [3:0] lut_324_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b0001011100011111;
    wire [3:0] lut_325_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b0100110100000000;
    wire [3:0] lut_326_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b1000101011101110;
    wire [3:0] lut_327_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b1100111100000100;
    wire [3:0] lut_328_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b0001011101111111;
    wire [3:0] lut_329_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b0100000011010101;
    wire [3:0] lut_330_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b0100110101010100;
    wire [3:0] lut_331_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b1110111010100000;
    wire [3:0] lut_332_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b1111111011101100;
    wire [3:0] lut_333_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b1101000011010101;
    wire [3:0] lut_334_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0001011101010111;
    wire [3:0] lut_335_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b0100010101000100;
    wire [3:0] lut_336_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b0001110100000010;
    wire [3:0] lut_337_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b1101111101000100;
    wire [3:0] lut_338_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b1110100011101010;
    wire [3:0] lut_339_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b1111000100010000;
    wire [3:0] lut_340_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b1110110011111110;
    wire [3:0] lut_341_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b0000000100001111;
    wire [3:0] lut_342_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b0001001100010001;
    wire [3:0] lut_343_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1111110011010100;
    wire [3:0] lut_344_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b0111000100010000;
    wire [3:0] lut_345_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b1110100011101100;
    wire [3:0] lut_346_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b0000001000101011;
    wire [3:0] lut_347_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0100110111111111;
    wire [3:0] lut_348_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b0000000100011111;
    wire [3:0] lut_349_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b1011001011110011;
    wire [3:0] lut_350_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b0001000000010001;
    wire [3:0] lut_351_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b0000010011001111;
    wire [3:0] lut_352_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b1010101110111111;
    wire [3:0] lut_353_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b0000000010101010;
    wire [3:0] lut_354_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b1010000010101000;
    wire [3:0] lut_355_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b0000000011001100;
    wire [3:0] lut_356_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b1110111010001110;
    wire [3:0] lut_357_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b1100110001000100;
    wire [3:0] lut_358_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b0000111110001111;
    wire [3:0] lut_359_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b0011111100001111;
    wire [3:0] lut_360_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b0010101000101011;
    wire [3:0] lut_361_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b0011011100111111;
    wire [3:0] lut_362_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b0111001100010001;
    wire [3:0] lut_363_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b0000000001011111;
    wire [3:0] lut_364_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b1110100010000000;
    wire [3:0] lut_365_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b1010101100101011;
    wire [3:0] lut_366_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b0101010001000000;
    wire [3:0] lut_367_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b1111000011110000;
    wire [3:0] lut_368_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b1100110101001101;
    wire [3:0] lut_369_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b1111000001110000;
    wire [3:0] lut_370_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b1010101011111111;
    wire [3:0] lut_371_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b0000010101011111;
    wire [3:0] lut_372_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b0101111101011111;
    wire [3:0] lut_373_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b0000000000101010;
    wire [3:0] lut_374_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b0001000111011111;
    wire [3:0] lut_375_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b0101010101110111;
    wire [3:0] lut_376_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b1111111100000111;
    wire [3:0] lut_377_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b0011001011110011;
    wire [3:0] lut_378_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1101010011111111;
    wire [3:0] lut_379_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b0011000001110001;
    wire [3:0] lut_380_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b0010101000101010;
    wire [3:0] lut_381_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b1000100011111010;
    wire [3:0] lut_382_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b1110111010000000;
    wire [3:0] lut_383_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0101110111011101;
    wire [3:0] lut_384_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b0100010101001101;
    wire [3:0] lut_385_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b0100111101001101;
    wire [3:0] lut_386_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b1011001111111111;
    wire [3:0] lut_387_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b1010101100100010;
    wire [3:0] lut_388_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b1010101011101010;
    wire [3:0] lut_389_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b0010001100100010;
    wire [3:0] lut_390_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b0000000011110100;
    wire [3:0] lut_391_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b1111001100110010;
    wire [3:0] lut_392_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b0011101100100010;
    wire [3:0] lut_393_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b0111011100010001;
    wire [3:0] lut_394_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b0011000001110011;
    wire [3:0] lut_395_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b0100111101001111;
    wire [3:0] lut_396_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b1000111100001010;
    wire [3:0] lut_397_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b1111111111111100;
    wire [3:0] lut_398_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b0000111100001100;
    wire [3:0] lut_399_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b0001000001110001;
    wire [3:0] lut_400_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b1010101011101110;
    wire [3:0] lut_401_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b0000111001001101;
    wire [3:0] lut_402_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b1111001111110001;
    wire [3:0] lut_403_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b0001111100000101;
    wire [3:0] lut_404_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b0000000100010111;
    wire [3:0] lut_405_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0111000111110011;
    wire [3:0] lut_406_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b1011001011111111;
    wire [3:0] lut_407_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b1010101000101010;
    wire [3:0] lut_408_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b1111101011101000;
    wire [3:0] lut_409_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b0111000111110101;
    wire [3:0] lut_410_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b0101011100010001;
    wire [3:0] lut_411_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b0010101100001010;
    wire [3:0] lut_412_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b1000110010001111;
    wire [3:0] lut_413_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0011011100000011;
    wire [3:0] lut_414_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b0100110101001100;
    wire [3:0] lut_415_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b0000010100010111;
    wire [3:0] lut_416_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b0001000011110001;
    wire [3:0] lut_417_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b0001011100010101;
    wire [3:0] lut_418_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b1111110101010000;
    wire [3:0] lut_419_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b0000000010111011;
    wire [3:0] lut_420_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b1011001110111011;
    wire [3:0] lut_421_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b1101010001010000;
    wire [3:0] lut_422_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b0001101100000000;
    wire [3:0] lut_423_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b0000011101111111;
    wire [3:0] lut_424_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b1011101100101010;
    wire [3:0] lut_425_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b0001010100000001;
    wire [3:0] lut_426_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b0001010100010111;
    wire [3:0] lut_427_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b0010111111111111;
    wire [3:0] lut_428_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b0000010001011111;
    wire [3:0] lut_429_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b0000011100111111;
    wire [3:0] lut_430_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b1111101000110010;
    wire [3:0] lut_431_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b0000111110111111;
    wire [3:0] lut_432_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b0100000011111100;
    wire [3:0] lut_433_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b1101010011110101;
    wire [3:0] lut_434_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b0011001100100011;
    wire [3:0] lut_435_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b1111001001100000;
    wire [3:0] lut_436_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b0001000100010111;
    wire [3:0] lut_437_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b1101010101000100;
    wire [3:0] lut_438_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b0011111100111111;
    wire [3:0] lut_439_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b1000111011101110;
    wire [3:0] lut_440_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b0000010001011111;
    wire [3:0] lut_441_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b1011101100100011;
    wire [3:0] lut_442_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1111001111111011;
    wire [3:0] lut_443_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b0011000101110111;
    wire [3:0] lut_444_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b1110111110001010;
    wire [3:0] lut_445_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b0010101100001010;
    wire [3:0] lut_446_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b1011101111110101;
    wire [3:0] lut_447_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b1111011100110001;
    wire [3:0] lut_448_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b1100110011011101;
    wire [3:0] lut_449_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b0010001100000010;
    wire [3:0] lut_450_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b0000000010001110;
    wire [3:0] lut_451_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b0100000001010000;
    wire [3:0] lut_452_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b1101110101010101;
    wire [3:0] lut_453_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0011000010110010;
    wire [3:0] lut_454_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b1010101011111011;
    wire [3:0] lut_455_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b0000000100010111;
    wire [3:0] lut_456_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b0000001010101011;
    wire [3:0] lut_457_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b0000100010101111;
    wire [3:0] lut_458_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b0101000111010111;
    wire [3:0] lut_459_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b0011000100010001;
    wire [3:0] lut_460_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b1111111111101000;
    wire [3:0] lut_461_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b0011001000111011;
    wire [3:0] lut_462_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b1011000100010000;
    wire [3:0] lut_463_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b1000101010001111;
    wire [3:0] lut_464_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b1111110011000000;
    wire [3:0] lut_465_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b1011011100101011;
    wire [3:0] lut_466_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1111110101000100;
    wire [3:0] lut_467_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b1000101010001011;
    wire [3:0] lut_468_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b0011001110110011;
    wire [3:0] lut_469_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b0000010100011111;
    wire [3:0] lut_470_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b1011101010100000;
    wire [3:0] lut_471_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b0000000011110011;
    wire [3:0] lut_472_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b0000001110111111;
    wire [3:0] lut_473_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b1100110110001000;
    wire [3:0] lut_474_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b1000111011101111;
    wire [3:0] lut_475_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b0011000000010001;
    wire [3:0] lut_476_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b1010111110001010;
    wire [3:0] lut_477_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b0011000011110011;
    wire [3:0] lut_478_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b1111111111111000;
    wire [3:0] lut_479_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b1000100010001100;
    wire [3:0] lut_480_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b1010101010101110;
    wire [3:0] lut_481_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b1101110001000100;
    wire [3:0] lut_482_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b1101000001010101;
    wire [3:0] lut_483_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b1101010001000000;
    wire [3:0] lut_484_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b0001011101011111;
    wire [3:0] lut_485_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b1111001011111111;
    wire [3:0] lut_486_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b0111001100010000;
    wire [3:0] lut_487_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1110111100001111;
    wire [3:0] lut_488_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b0101011101011111;
    wire [3:0] lut_489_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b0100010011010100;
    wire [3:0] lut_490_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b0010001010101011;
    wire [3:0] lut_491_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b1000111100001111;
    wire [3:0] lut_492_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b0000000100010111;
    wire [3:0] lut_493_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b0111000011110001;
    wire [3:0] lut_494_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b1100100011001000;
    wire [3:0] lut_495_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b1101010101000000;
    wire [3:0] lut_496_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b0000111000001110;
    wire [3:0] lut_497_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b0101110101001101;
    wire [3:0] lut_498_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b1110100011111110;
    wire [3:0] lut_499_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b0111011101110111;
    wire [3:0] lut_500_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b1101011100000000;
    wire [3:0] lut_501_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b1111010111110000;
    wire [3:0] lut_502_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b0000110011101111;
    wire [3:0] lut_503_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b1111110111110100;
    wire [3:0] lut_504_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b0111000000010000;
    wire [3:0] lut_505_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b1100010011111100;
    wire [3:0] lut_506_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b1111101100100000;
    wire [3:0] lut_507_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b0011001000100000;
    wire [3:0] lut_508_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b1111111011001100;
    wire [3:0] lut_509_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b0010101110111011;
    wire [3:0] lut_510_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0000001100111011;
    wire [3:0] lut_511_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [15:0] lut_512_table = 16'b1111101000110000;
    wire [3:0] lut_512_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [15:0] lut_513_table = 16'b0011101100111011;
    wire [3:0] lut_513_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [15:0] lut_514_table = 16'b1111010111110011;
    wire [3:0] lut_514_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [15:0] lut_515_table = 16'b1010000011110000;
    wire [3:0] lut_515_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [15:0] lut_516_table = 16'b0010101100001111;
    wire [3:0] lut_516_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [15:0] lut_517_table = 16'b0101000101110001;
    wire [3:0] lut_517_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [15:0] lut_518_table = 16'b0010001011111011;
    wire [3:0] lut_518_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [15:0] lut_519_table = 16'b0010001000101010;
    wire [3:0] lut_519_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [15:0] lut_520_table = 16'b0010001100000011;
    wire [3:0] lut_520_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [15:0] lut_521_table = 16'b0000100010001111;
    wire [3:0] lut_521_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [15:0] lut_522_table = 16'b1110100001000000;
    wire [3:0] lut_522_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [15:0] lut_523_table = 16'b0000110010101110;
    wire [3:0] lut_523_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [15:0] lut_524_table = 16'b0000000001011111;
    wire [3:0] lut_524_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [15:0] lut_525_table = 16'b0001011111111111;
    wire [3:0] lut_525_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [15:0] lut_526_table = 16'b0111010001110101;
    wire [3:0] lut_526_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [15:0] lut_527_table = 16'b0101010100000000;
    wire [3:0] lut_527_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [15:0] lut_528_table = 16'b1111000011110000;
    wire [3:0] lut_528_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [15:0] lut_529_table = 16'b1101010011010101;
    wire [3:0] lut_529_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [15:0] lut_530_table = 16'b0000111011001111;
    wire [3:0] lut_530_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [15:0] lut_531_table = 16'b1010101010111111;
    wire [3:0] lut_531_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [15:0] lut_532_table = 16'b0100010111010111;
    wire [3:0] lut_532_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [15:0] lut_533_table = 16'b1110111100000000;
    wire [3:0] lut_533_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [15:0] lut_534_table = 16'b0000000010101010;
    wire [3:0] lut_534_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [15:0] lut_535_table = 16'b1010101010101000;
    wire [3:0] lut_535_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [15:0] lut_536_table = 16'b1111100000000000;
    wire [3:0] lut_536_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [15:0] lut_537_table = 16'b1000000011111010;
    wire [3:0] lut_537_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [15:0] lut_538_table = 16'b0000101010101110;
    wire [3:0] lut_538_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [15:0] lut_539_table = 16'b0100010100000000;
    wire [3:0] lut_539_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [15:0] lut_540_table = 16'b0000000011110101;
    wire [3:0] lut_540_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [15:0] lut_541_table = 16'b1000001010111011;
    wire [3:0] lut_541_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [15:0] lut_542_table = 16'b1000000011111110;
    wire [3:0] lut_542_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [15:0] lut_543_table = 16'b1110100011000000;
    wire [3:0] lut_543_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [15:0] lut_544_table = 16'b0100110111111111;
    wire [3:0] lut_544_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [15:0] lut_545_table = 16'b1011001010111011;
    wire [3:0] lut_545_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [15:0] lut_546_table = 16'b0010000000110011;
    wire [3:0] lut_546_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [15:0] lut_547_table = 16'b0100110100000100;
    wire [3:0] lut_547_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [15:0] lut_548_table = 16'b0000101100101011;
    wire [3:0] lut_548_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [15:0] lut_549_table = 16'b0011111101111111;
    wire [3:0] lut_549_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [15:0] lut_550_table = 16'b0100110111011101;
    wire [3:0] lut_550_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [15:0] lut_551_table = 16'b1011111100001111;
    wire [3:0] lut_551_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [15:0] lut_552_table = 16'b0000110011001101;
    wire [3:0] lut_552_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [15:0] lut_553_table = 16'b0011111100110011;
    wire [3:0] lut_553_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [15:0] lut_554_table = 16'b1000100010101110;
    wire [3:0] lut_554_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [15:0] lut_555_table = 16'b0010001010111011;
    wire [3:0] lut_555_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [15:0] lut_556_table = 16'b1011001000100000;
    wire [3:0] lut_556_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [15:0] lut_557_table = 16'b1000111100001010;
    wire [3:0] lut_557_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [15:0] lut_558_table = 16'b0000001000101010;
    wire [3:0] lut_558_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [15:0] lut_559_table = 16'b1110110011111111;
    wire [3:0] lut_559_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [15:0] lut_560_table = 16'b0100000011110111;
    wire [3:0] lut_560_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [15:0] lut_561_table = 16'b1100010011000100;
    wire [3:0] lut_561_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [15:0] lut_562_table = 16'b1011111100101011;
    wire [3:0] lut_562_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [15:0] lut_563_table = 16'b0000000011101100;
    wire [3:0] lut_563_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [15:0] lut_564_table = 16'b0011101000000010;
    wire [3:0] lut_564_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [15:0] lut_565_table = 16'b0000000100010111;
    wire [3:0] lut_565_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [15:0] lut_566_table = 16'b0010101010111111;
    wire [3:0] lut_566_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [15:0] lut_567_table = 16'b0101010101010100;
    wire [3:0] lut_567_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [15:0] lut_568_table = 16'b0010000010110011;
    wire [3:0] lut_568_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [15:0] lut_569_table = 16'b1111101011101000;
    wire [3:0] lut_569_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [15:0] lut_570_table = 16'b0001001111110111;
    wire [3:0] lut_570_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [15:0] lut_571_table = 16'b1100000011101100;
    wire [3:0] lut_571_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [15:0] lut_572_table = 16'b0111000011110111;
    wire [3:0] lut_572_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [15:0] lut_573_table = 16'b1000110010001111;
    wire [3:0] lut_573_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [15:0] lut_574_table = 16'b1110111010000000;
    wire [3:0] lut_574_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [15:0] lut_575_table = 16'b1011000010111011;
    wire [3:0] lut_575_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [15:0] lut_576_table = 16'b1111101011111000;
    wire [3:0] lut_576_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [15:0] lut_577_table = 16'b1010100011111011;
    wire [3:0] lut_577_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [15:0] lut_578_table = 16'b1110100011101000;
    wire [3:0] lut_578_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [15:0] lut_579_table = 16'b1100110011111111;
    wire [3:0] lut_579_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [15:0] lut_580_table = 16'b0000111100001011;
    wire [3:0] lut_580_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [15:0] lut_581_table = 16'b0011001110110011;
    wire [3:0] lut_581_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [15:0] lut_582_table = 16'b0010001000111011;
    wire [3:0] lut_582_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [15:0] lut_583_table = 16'b1000100011101100;
    wire [3:0] lut_583_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [15:0] lut_584_table = 16'b1111101010000000;
    wire [3:0] lut_584_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [15:0] lut_585_table = 16'b0010001011111010;
    wire [3:0] lut_585_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [15:0] lut_586_table = 16'b1110100011111110;
    wire [3:0] lut_586_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [15:0] lut_587_table = 16'b0001011101010111;
    wire [3:0] lut_587_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [15:0] lut_588_table = 16'b0010101111111111;
    wire [3:0] lut_588_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [15:0] lut_589_table = 16'b0000001100010111;
    wire [3:0] lut_589_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [15:0] lut_590_table = 16'b1111111010000000;
    wire [3:0] lut_590_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [15:0] lut_591_table = 16'b1111111111110000;
    wire [3:0] lut_591_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [15:0] lut_592_table = 16'b1011001110110010;
    wire [3:0] lut_592_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [15:0] lut_593_table = 16'b1010111000001010;
    wire [3:0] lut_593_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [15:0] lut_594_table = 16'b0000000011001100;
    wire [3:0] lut_594_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [15:0] lut_595_table = 16'b0111000111110101;
    wire [3:0] lut_595_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [15:0] lut_596_table = 16'b0000010100010101;
    wire [3:0] lut_596_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [15:0] lut_597_table = 16'b0001011100110111;
    wire [3:0] lut_597_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [15:0] lut_598_table = 16'b1101010100000000;
    wire [3:0] lut_598_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [15:0] lut_599_table = 16'b1011101110101010;
    wire [3:0] lut_599_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [15:0] lut_600_table = 16'b1000111011101111;
    wire [3:0] lut_600_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [15:0] lut_601_table = 16'b1111101110100000;
    wire [3:0] lut_601_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [15:0] lut_602_table = 16'b1100000011000000;
    wire [3:0] lut_602_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [15:0] lut_603_table = 16'b1011000011111011;
    wire [3:0] lut_603_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [15:0] lut_604_table = 16'b0011000011110111;
    wire [3:0] lut_604_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [15:0] lut_605_table = 16'b1111111110001010;
    wire [3:0] lut_605_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [15:0] lut_606_table = 16'b1111010100110011;
    wire [3:0] lut_606_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [15:0] lut_607_table = 16'b1111010101010000;
    wire [3:0] lut_607_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [15:0] lut_608_table = 16'b0000111011001110;
    wire [3:0] lut_608_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [15:0] lut_609_table = 16'b1101111100001101;
    wire [3:0] lut_609_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [15:0] lut_610_table = 16'b0101010111110111;
    wire [3:0] lut_610_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [15:0] lut_611_table = 16'b0000000000001110;
    wire [3:0] lut_611_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [15:0] lut_612_table = 16'b0000110011011111;
    wire [3:0] lut_612_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [15:0] lut_613_table = 16'b0110000011101010;
    wire [3:0] lut_613_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [15:0] lut_614_table = 16'b0011000000110010;
    wire [3:0] lut_614_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [15:0] lut_615_table = 16'b1101110001000100;
    wire [3:0] lut_615_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [15:0] lut_616_table = 16'b0000000100010111;
    wire [3:0] lut_616_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [15:0] lut_617_table = 16'b1111110111110100;
    wire [3:0] lut_617_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [15:0] lut_618_table = 16'b0101010101110111;
    wire [3:0] lut_618_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [15:0] lut_619_table = 16'b1010101010101010;
    wire [3:0] lut_619_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [15:0] lut_620_table = 16'b0111001000000000;
    wire [3:0] lut_620_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [15:0] lut_621_table = 16'b0000001100000011;
    wire [3:0] lut_621_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [15:0] lut_622_table = 16'b0011001100110010;
    wire [3:0] lut_622_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [15:0] lut_623_table = 16'b1100110011101111;
    wire [3:0] lut_623_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [15:0] lut_624_table = 16'b1111011101110101;
    wire [3:0] lut_624_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [15:0] lut_625_table = 16'b1111110011000000;
    wire [3:0] lut_625_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [15:0] lut_626_table = 16'b0001000011110011;
    wire [3:0] lut_626_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [15:0] lut_627_table = 16'b0000001000111111;
    wire [3:0] lut_627_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [15:0] lut_628_table = 16'b0011000001110000;
    wire [3:0] lut_628_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [15:0] lut_629_table = 16'b1010111100000001;
    wire [3:0] lut_629_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [15:0] lut_630_table = 16'b1000100011101110;
    wire [3:0] lut_630_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [15:0] lut_631_table = 16'b1011000000100000;
    wire [3:0] lut_631_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [15:0] lut_632_table = 16'b0001010101111111;
    wire [3:0] lut_632_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [15:0] lut_633_table = 16'b1111010011010000;
    wire [3:0] lut_633_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [15:0] lut_634_table = 16'b0000010101010101;
    wire [3:0] lut_634_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [15:0] lut_635_table = 16'b0111001100110000;
    wire [3:0] lut_635_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [15:0] lut_636_table = 16'b1110111110001110;
    wire [3:0] lut_636_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [15:0] lut_637_table = 16'b0101000001110101;
    wire [3:0] lut_637_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [15:0] lut_638_table = 16'b1010101000100010;
    wire [3:0] lut_638_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [15:0] lut_639_table = 16'b0001000100010111;
    wire [3:0] lut_639_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub5
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        639:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        639:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub5_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub5_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub5_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [639:0]  in_data,
            output wire [639:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1011001010110010;
    wire [3:0] lut_0_select = {
                             in_data[459],
                             in_data[432],
                             in_data[227],
                             in_data[285]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b0000001011111111;
    wire [3:0] lut_1_select = {
                             in_data[4],
                             in_data[246],
                             in_data[502],
                             in_data[312]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b1111101011111010;
    wire [3:0] lut_2_select = {
                             in_data[638],
                             in_data[287],
                             in_data[633],
                             in_data[148]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1100110011111111;
    wire [3:0] lut_3_select = {
                             in_data[507],
                             in_data[175],
                             in_data[521],
                             in_data[590]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b1110111010000100;
    wire [3:0] lut_4_select = {
                             in_data[413],
                             in_data[153],
                             in_data[196],
                             in_data[123]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b0000001100101111;
    wire [3:0] lut_5_select = {
                             in_data[99],
                             in_data[212],
                             in_data[608],
                             in_data[105]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b1010111100000111;
    wire [3:0] lut_6_select = {
                             in_data[71],
                             in_data[252],
                             in_data[98],
                             in_data[551]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b0011111100000000;
    wire [3:0] lut_7_select = {
                             in_data[357],
                             in_data[43],
                             in_data[419],
                             in_data[199]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1111000001000000;
    wire [3:0] lut_8_select = {
                             in_data[606],
                             in_data[247],
                             in_data[472],
                             in_data[19]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b1100000011000000;
    wire [3:0] lut_9_select = {
                             in_data[211],
                             in_data[586],
                             in_data[163],
                             in_data[433]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b1101010011010101;
    wire [3:0] lut_10_select = {
                             in_data[569],
                             in_data[381],
                             in_data[441],
                             in_data[429]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b1101000011110000;
    wire [3:0] lut_11_select = {
                             in_data[282],
                             in_data[438],
                             in_data[360],
                             in_data[113]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b0000110011001100;
    wire [3:0] lut_12_select = {
                             in_data[207],
                             in_data[451],
                             in_data[359],
                             in_data[585]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0000000000000101;
    wire [3:0] lut_13_select = {
                             in_data[155],
                             in_data[293],
                             in_data[573],
                             in_data[42]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0100010011010100;
    wire [3:0] lut_14_select = {
                             in_data[25],
                             in_data[146],
                             in_data[292],
                             in_data[192]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1101110100000000;
    wire [3:0] lut_15_select = {
                             in_data[92],
                             in_data[388],
                             in_data[603],
                             in_data[430]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b0000101100110011;
    wire [3:0] lut_16_select = {
                             in_data[93],
                             in_data[575],
                             in_data[464],
                             in_data[232]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b0111111101010101;
    wire [3:0] lut_17_select = {
                             in_data[520],
                             in_data[300],
                             in_data[107],
                             in_data[504]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0001000100000001;
    wire [3:0] lut_18_select = {
                             in_data[242],
                             in_data[161],
                             in_data[533],
                             in_data[324]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b1100110010001100;
    wire [3:0] lut_19_select = {
                             in_data[129],
                             in_data[594],
                             in_data[330],
                             in_data[114]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0000110100001111;
    wire [3:0] lut_20_select = {
                             in_data[144],
                             in_data[637],
                             in_data[343],
                             in_data[183]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b1111111100101011;
    wire [3:0] lut_21_select = {
                             in_data[185],
                             in_data[191],
                             in_data[170],
                             in_data[208]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b1011001111110011;
    wire [3:0] lut_22_select = {
                             in_data[344],
                             in_data[220],
                             in_data[371],
                             in_data[261]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0101110101010100;
    wire [3:0] lut_23_select = {
                             in_data[409],
                             in_data[178],
                             in_data[281],
                             in_data[498]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1011101110111011;
    wire [3:0] lut_24_select = {
                             in_data[34],
                             in_data[122],
                             in_data[214],
                             in_data[505]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0001010101110001;
    wire [3:0] lut_25_select = {
                             in_data[296],
                             in_data[591],
                             in_data[598],
                             in_data[424]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b0010001010101010;
    wire [3:0] lut_26_select = {
                             in_data[313],
                             in_data[154],
                             in_data[530],
                             in_data[570]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1111111010001000;
    wire [3:0] lut_27_select = {
                             in_data[222],
                             in_data[609],
                             in_data[280],
                             in_data[66]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b0000111010001110;
    wire [3:0] lut_28_select = {
                             in_data[83],
                             in_data[494],
                             in_data[140],
                             in_data[69]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b1100110100000100;
    wire [3:0] lut_29_select = {
                             in_data[37],
                             in_data[180],
                             in_data[600],
                             in_data[532]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b1000100010001000;
    wire [3:0] lut_30_select = {
                             in_data[40],
                             in_data[514],
                             in_data[64],
                             in_data[453]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1101111111011100;
    wire [3:0] lut_31_select = {
                             in_data[310],
                             in_data[230],
                             in_data[528],
                             in_data[455]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b1010101010101010;
    wire [3:0] lut_32_select = {
                             in_data[583],
                             in_data[260],
                             in_data[560],
                             in_data[412]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b0101110101000101;
    wire [3:0] lut_33_select = {
                             in_data[24],
                             in_data[461],
                             in_data[68],
                             in_data[82]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1111001110110011;
    wire [3:0] lut_34_select = {
                             in_data[350],
                             in_data[307],
                             in_data[120],
                             in_data[20]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b0100111111001100;
    wire [3:0] lut_35_select = {
                             in_data[554],
                             in_data[632],
                             in_data[595],
                             in_data[563]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b1101010011010100;
    wire [3:0] lut_36_select = {
                             in_data[431],
                             in_data[386],
                             in_data[354],
                             in_data[164]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0101010111010100;
    wire [3:0] lut_37_select = {
                             in_data[284],
                             in_data[512],
                             in_data[139],
                             in_data[26]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b0000000111111111;
    wire [3:0] lut_38_select = {
                             in_data[204],
                             in_data[380],
                             in_data[465],
                             in_data[210]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0101000111111111;
    wire [3:0] lut_39_select = {
                             in_data[397],
                             in_data[390],
                             in_data[97],
                             in_data[221]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b1011111100000011;
    wire [3:0] lut_40_select = {
                             in_data[198],
                             in_data[500],
                             in_data[104],
                             in_data[422]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b1011001100100010;
    wire [3:0] lut_41_select = {
                             in_data[151],
                             in_data[63],
                             in_data[538],
                             in_data[111]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b1101110111011101;
    wire [3:0] lut_42_select = {
                             in_data[336],
                             in_data[171],
                             in_data[395],
                             in_data[270]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0000110001001100;
    wire [3:0] lut_43_select = {
                             in_data[11],
                             in_data[169],
                             in_data[301],
                             in_data[394]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b0100110011001100;
    wire [3:0] lut_44_select = {
                             in_data[50],
                             in_data[478],
                             in_data[233],
                             in_data[264]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b1100111100010101;
    wire [3:0] lut_45_select = {
                             in_data[238],
                             in_data[321],
                             in_data[138],
                             in_data[486]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b0100110011001100;
    wire [3:0] lut_46_select = {
                             in_data[450],
                             in_data[434],
                             in_data[517],
                             in_data[546]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b0001011100010111;
    wire [3:0] lut_47_select = {
                             in_data[9],
                             in_data[1],
                             in_data[383],
                             in_data[278]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b1111111101000100;
    wire [3:0] lut_48_select = {
                             in_data[224],
                             in_data[249],
                             in_data[414],
                             in_data[579]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b1010101000100000;
    wire [3:0] lut_49_select = {
                             in_data[187],
                             in_data[543],
                             in_data[124],
                             in_data[541]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0101111100000111;
    wire [3:0] lut_50_select = {
                             in_data[518],
                             in_data[197],
                             in_data[471],
                             in_data[561]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b0000001001111111;
    wire [3:0] lut_51_select = {
                             in_data[240],
                             in_data[589],
                             in_data[635],
                             in_data[341]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1111111100110000;
    wire [3:0] lut_52_select = {
                             in_data[411],
                             in_data[30],
                             in_data[447],
                             in_data[339]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b0101000100010000;
    wire [3:0] lut_53_select = {
                             in_data[477],
                             in_data[147],
                             in_data[338],
                             in_data[62]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b0101111100001101;
    wire [3:0] lut_54_select = {
                             in_data[580],
                             in_data[346],
                             in_data[168],
                             in_data[203]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b1111110111010100;
    wire [3:0] lut_55_select = {
                             in_data[558],
                             in_data[226],
                             in_data[487],
                             in_data[488]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b1111000000010000;
    wire [3:0] lut_56_select = {
                             in_data[5],
                             in_data[298],
                             in_data[127],
                             in_data[476]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b1000000010101010;
    wire [3:0] lut_57_select = {
                             in_data[454],
                             in_data[315],
                             in_data[448],
                             in_data[27]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b1111101010111000;
    wire [3:0] lut_58_select = {
                             in_data[463],
                             in_data[65],
                             in_data[536],
                             in_data[255]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b0000000011111110;
    wire [3:0] lut_59_select = {
                             in_data[160],
                             in_data[45],
                             in_data[392],
                             in_data[539]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b1000111010101000;
    wire [3:0] lut_60_select = {
                             in_data[28],
                             in_data[391],
                             in_data[529],
                             in_data[218]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b1011101000100010;
    wire [3:0] lut_61_select = {
                             in_data[345],
                             in_data[581],
                             in_data[557],
                             in_data[481]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b1000100010001000;
    wire [3:0] lut_62_select = {
                             in_data[480],
                             in_data[425],
                             in_data[250],
                             in_data[396]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b1010101010001000;
    wire [3:0] lut_63_select = {
                             in_data[248],
                             in_data[58],
                             in_data[545],
                             in_data[624]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b1111101000100000;
    wire [3:0] lut_64_select = {
                             in_data[70],
                             in_data[88],
                             in_data[442],
                             in_data[439]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b1010101010101010;
    wire [3:0] lut_65_select = {
                             in_data[437],
                             in_data[95],
                             in_data[17],
                             in_data[382]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b1010111110001111;
    wire [3:0] lut_66_select = {
                             in_data[564],
                             in_data[179],
                             in_data[121],
                             in_data[510]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b1101010101000100;
    wire [3:0] lut_67_select = {
                             in_data[7],
                             in_data[59],
                             in_data[332],
                             in_data[374]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b1110110011101000;
    wire [3:0] lut_68_select = {
                             in_data[491],
                             in_data[402],
                             in_data[616],
                             in_data[614]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b0011000011110011;
    wire [3:0] lut_69_select = {
                             in_data[254],
                             in_data[209],
                             in_data[446],
                             in_data[239]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b1010101110111011;
    wire [3:0] lut_70_select = {
                             in_data[599],
                             in_data[256],
                             in_data[231],
                             in_data[547]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0111011000010000;
    wire [3:0] lut_71_select = {
                             in_data[612],
                             in_data[152],
                             in_data[410],
                             in_data[368]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b1010101010101010;
    wire [3:0] lut_72_select = {
                             in_data[131],
                             in_data[143],
                             in_data[316],
                             in_data[35]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b0000111010101111;
    wire [3:0] lut_73_select = {
                             in_data[277],
                             in_data[13],
                             in_data[337],
                             in_data[184]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0001001100110011;
    wire [3:0] lut_74_select = {
                             in_data[400],
                             in_data[12],
                             in_data[605],
                             in_data[349]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b1101000011111000;
    wire [3:0] lut_75_select = {
                             in_data[23],
                             in_data[362],
                             in_data[162],
                             in_data[537]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0001000011111101;
    wire [3:0] lut_76_select = {
                             in_data[376],
                             in_data[94],
                             in_data[331],
                             in_data[492]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b0000001100000011;
    wire [3:0] lut_77_select = {
                             in_data[286],
                             in_data[55],
                             in_data[358],
                             in_data[257]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b1111101010001000;
    wire [3:0] lut_78_select = {
                             in_data[513],
                             in_data[39],
                             in_data[617],
                             in_data[565]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b1111001110110000;
    wire [3:0] lut_79_select = {
                             in_data[577],
                             in_data[290],
                             in_data[452],
                             in_data[630]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b1100111010001100;
    wire [3:0] lut_80_select = {
                             in_data[615],
                             in_data[87],
                             in_data[351],
                             in_data[302]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b1111010101010000;
    wire [3:0] lut_81_select = {
                             in_data[370],
                             in_data[550],
                             in_data[172],
                             in_data[493]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1111000011110000;
    wire [3:0] lut_82_select = {
                             in_data[456],
                             in_data[108],
                             in_data[317],
                             in_data[84]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b1101010101010101;
    wire [3:0] lut_83_select = {
                             in_data[291],
                             in_data[258],
                             in_data[613],
                             in_data[320]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b1111111110100000;
    wire [3:0] lut_84_select = {
                             in_data[323],
                             in_data[484],
                             in_data[259],
                             in_data[289]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b0111010101110110;
    wire [3:0] lut_85_select = {
                             in_data[311],
                             in_data[629],
                             in_data[523],
                             in_data[457]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b0010101100111011;
    wire [3:0] lut_86_select = {
                             in_data[469],
                             in_data[496],
                             in_data[335],
                             in_data[333]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b1110000011100000;
    wire [3:0] lut_87_select = {
                             in_data[596],
                             in_data[375],
                             in_data[398],
                             in_data[318]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b0111010101010001;
    wire [3:0] lut_88_select = {
                             in_data[135],
                             in_data[253],
                             in_data[423],
                             in_data[475]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b1101010101000000;
    wire [3:0] lut_89_select = {
                             in_data[283],
                             in_data[117],
                             in_data[265],
                             in_data[623]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b1111101011111010;
    wire [3:0] lut_90_select = {
                             in_data[126],
                             in_data[522],
                             in_data[156],
                             in_data[445]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b1111001010110000;
    wire [3:0] lut_91_select = {
                             in_data[200],
                             in_data[406],
                             in_data[194],
                             in_data[468]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b1110100010101000;
    wire [3:0] lut_92_select = {
                             in_data[201],
                             in_data[149],
                             in_data[219],
                             in_data[404]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0010101110101011;
    wire [3:0] lut_93_select = {
                             in_data[96],
                             in_data[567],
                             in_data[15],
                             in_data[6]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b0000001100000011;
    wire [3:0] lut_94_select = {
                             in_data[150],
                             in_data[552],
                             in_data[625],
                             in_data[263]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b1110010011100100;
    wire [3:0] lut_95_select = {
                             in_data[85],
                             in_data[458],
                             in_data[542],
                             in_data[553]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1111111010000000;
    wire [3:0] lut_96_select = {
                             in_data[426],
                             in_data[319],
                             in_data[89],
                             in_data[288]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b0000110100001101;
    wire [3:0] lut_97_select = {
                             in_data[473],
                             in_data[444],
                             in_data[91],
                             in_data[628]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1111001101110001;
    wire [3:0] lut_98_select = {
                             in_data[262],
                             in_data[166],
                             in_data[495],
                             in_data[639]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b1000110000001000;
    wire [3:0] lut_99_select = {
                             in_data[408],
                             in_data[101],
                             in_data[379],
                             in_data[141]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b1000111011001111;
    wire [3:0] lut_100_select = {
                             in_data[32],
                             in_data[571],
                             in_data[145],
                             in_data[49]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b1100110001001100;
    wire [3:0] lut_101_select = {
                             in_data[0],
                             in_data[470],
                             in_data[420],
                             in_data[627]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b0000001100100111;
    wire [3:0] lut_102_select = {
                             in_data[213],
                             in_data[393],
                             in_data[86],
                             in_data[142]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1111001010110000;
    wire [3:0] lut_103_select = {
                             in_data[77],
                             in_data[369],
                             in_data[556],
                             in_data[416]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b0100010001001101;
    wire [3:0] lut_104_select = {
                             in_data[622],
                             in_data[314],
                             in_data[237],
                             in_data[356]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1101010011010000;
    wire [3:0] lut_105_select = {
                             in_data[509],
                             in_data[190],
                             in_data[167],
                             in_data[544]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b1111000011111110;
    wire [3:0] lut_106_select = {
                             in_data[578],
                             in_data[340],
                             in_data[462],
                             in_data[427]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b1111000011111111;
    wire [3:0] lut_107_select = {
                             in_data[322],
                             in_data[587],
                             in_data[8],
                             in_data[159]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b0111000001010101;
    wire [3:0] lut_108_select = {
                             in_data[515],
                             in_data[574],
                             in_data[325],
                             in_data[519]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b1011000011111010;
    wire [3:0] lut_109_select = {
                             in_data[436],
                             in_data[125],
                             in_data[593],
                             in_data[29]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b0000011101111111;
    wire [3:0] lut_110_select = {
                             in_data[112],
                             in_data[56],
                             in_data[53],
                             in_data[72]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000101100001111;
    wire [3:0] lut_111_select = {
                             in_data[631],
                             in_data[132],
                             in_data[46],
                             in_data[118]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b1011000011110000;
    wire [3:0] lut_112_select = {
                             in_data[243],
                             in_data[216],
                             in_data[276],
                             in_data[206]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b0000011101111111;
    wire [3:0] lut_113_select = {
                             in_data[116],
                             in_data[449],
                             in_data[54],
                             in_data[103]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1000111010111100;
    wire [3:0] lut_114_select = {
                             in_data[610],
                             in_data[14],
                             in_data[361],
                             in_data[274]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0000001010101011;
    wire [3:0] lut_115_select = {
                             in_data[269],
                             in_data[205],
                             in_data[267],
                             in_data[562]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b1111111111110000;
    wire [3:0] lut_116_select = {
                             in_data[548],
                             in_data[268],
                             in_data[531],
                             in_data[372]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b1100000011111101;
    wire [3:0] lut_117_select = {
                             in_data[499],
                             in_data[225],
                             in_data[634],
                             in_data[67]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1111100010000000;
    wire [3:0] lut_118_select = {
                             in_data[158],
                             in_data[173],
                             in_data[294],
                             in_data[78]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b1010101010110010;
    wire [3:0] lut_119_select = {
                             in_data[328],
                             in_data[421],
                             in_data[527],
                             in_data[90]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b1010000010100000;
    wire [3:0] lut_120_select = {
                             in_data[621],
                             in_data[309],
                             in_data[130],
                             in_data[348]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b0000011100000111;
    wire [3:0] lut_121_select = {
                             in_data[186],
                             in_data[460],
                             in_data[182],
                             in_data[607]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b0000101100011111;
    wire [3:0] lut_122_select = {
                             in_data[566],
                             in_data[48],
                             in_data[308],
                             in_data[241]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b0000111110101111;
    wire [3:0] lut_123_select = {
                             in_data[51],
                             in_data[272],
                             in_data[501],
                             in_data[474]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b0000001010111111;
    wire [3:0] lut_124_select = {
                             in_data[251],
                             in_data[188],
                             in_data[385],
                             in_data[52]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b1011001010110010;
    wire [3:0] lut_125_select = {
                             in_data[636],
                             in_data[535],
                             in_data[2],
                             in_data[195]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b0101010111110101;
    wire [3:0] lut_126_select = {
                             in_data[100],
                             in_data[244],
                             in_data[279],
                             in_data[326]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0000000001110101;
    wire [3:0] lut_127_select = {
                             in_data[177],
                             in_data[18],
                             in_data[355],
                             in_data[597]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b1000110001001111;
    wire [3:0] lut_128_select = {
                             in_data[271],
                             in_data[582],
                             in_data[128],
                             in_data[295]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b0000100010101111;
    wire [3:0] lut_129_select = {
                             in_data[619],
                             in_data[215],
                             in_data[626],
                             in_data[568]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b1111111110110010;
    wire [3:0] lut_130_select = {
                             in_data[57],
                             in_data[378],
                             in_data[329],
                             in_data[347]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b1010111110000000;
    wire [3:0] lut_131_select = {
                             in_data[364],
                             in_data[10],
                             in_data[31],
                             in_data[235]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b1100110011111111;
    wire [3:0] lut_132_select = {
                             in_data[106],
                             in_data[136],
                             in_data[466],
                             in_data[440]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0101010101010101;
    wire [3:0] lut_133_select = {
                             in_data[373],
                             in_data[110],
                             in_data[176],
                             in_data[482]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b0001010100010001;
    wire [3:0] lut_134_select = {
                             in_data[584],
                             in_data[479],
                             in_data[490],
                             in_data[181]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b1011111100100011;
    wire [3:0] lut_135_select = {
                             in_data[485],
                             in_data[559],
                             in_data[428],
                             in_data[102]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b1111111111001100;
    wire [3:0] lut_136_select = {
                             in_data[299],
                             in_data[119],
                             in_data[229],
                             in_data[503]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b0101000011110011;
    wire [3:0] lut_137_select = {
                             in_data[525],
                             in_data[327],
                             in_data[61],
                             in_data[60]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b0010101100100011;
    wire [3:0] lut_138_select = {
                             in_data[76],
                             in_data[511],
                             in_data[534],
                             in_data[75]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b0000010111111111;
    wire [3:0] lut_139_select = {
                             in_data[189],
                             in_data[506],
                             in_data[266],
                             in_data[137]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b1010101011111011;
    wire [3:0] lut_140_select = {
                             in_data[47],
                             in_data[16],
                             in_data[41],
                             in_data[497]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b1000101001001110;
    wire [3:0] lut_141_select = {
                             in_data[236],
                             in_data[601],
                             in_data[303],
                             in_data[443]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b1111000011111100;
    wire [3:0] lut_142_select = {
                             in_data[273],
                             in_data[38],
                             in_data[165],
                             in_data[555]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0010000011110000;
    wire [3:0] lut_143_select = {
                             in_data[611],
                             in_data[592],
                             in_data[304],
                             in_data[352]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b1101110101000000;
    wire [3:0] lut_144_select = {
                             in_data[157],
                             in_data[618],
                             in_data[403],
                             in_data[228]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b1011111110001000;
    wire [3:0] lut_145_select = {
                             in_data[44],
                             in_data[3],
                             in_data[405],
                             in_data[387]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1111001110100010;
    wire [3:0] lut_146_select = {
                             in_data[526],
                             in_data[245],
                             in_data[234],
                             in_data[483]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0010101100100011;
    wire [3:0] lut_147_select = {
                             in_data[133],
                             in_data[367],
                             in_data[115],
                             in_data[22]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b1010001011111111;
    wire [3:0] lut_148_select = {
                             in_data[275],
                             in_data[81],
                             in_data[79],
                             in_data[365]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b1111001100110000;
    wire [3:0] lut_149_select = {
                             in_data[417],
                             in_data[353],
                             in_data[134],
                             in_data[174]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b1010101010111010;
    wire [3:0] lut_150_select = {
                             in_data[202],
                             in_data[36],
                             in_data[572],
                             in_data[604]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b0010000011110011;
    wire [3:0] lut_151_select = {
                             in_data[549],
                             in_data[389],
                             in_data[588],
                             in_data[407]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b0011001011111111;
    wire [3:0] lut_152_select = {
                             in_data[489],
                             in_data[576],
                             in_data[540],
                             in_data[297]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1000100011111010;
    wire [3:0] lut_153_select = {
                             in_data[342],
                             in_data[602],
                             in_data[384],
                             in_data[21]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0000111100001111;
    wire [3:0] lut_154_select = {
                             in_data[193],
                             in_data[377],
                             in_data[415],
                             in_data[109]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b1111101011111000;
    wire [3:0] lut_155_select = {
                             in_data[418],
                             in_data[516],
                             in_data[366],
                             in_data[217]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b1101110101000100;
    wire [3:0] lut_156_select = {
                             in_data[620],
                             in_data[399],
                             in_data[435],
                             in_data[305]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b0010000010110010;
    wire [3:0] lut_157_select = {
                             in_data[508],
                             in_data[524],
                             in_data[334],
                             in_data[401]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b0000000011110101;
    wire [3:0] lut_158_select = {
                             in_data[467],
                             in_data[223],
                             in_data[80],
                             in_data[74]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b0000001100010011;
    wire [3:0] lut_159_select = {
                             in_data[33],
                             in_data[73],
                             in_data[363],
                             in_data[306]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
    
    // LUT : 160
    wire [15:0] lut_160_table = 16'b1101111101011101;
    wire [3:0] lut_160_select = {
                             in_data[303],
                             in_data[411],
                             in_data[252],
                             in_data[325]};
    
    wire lut_160_out = lut_160_table[lut_160_select];
    
    generate
    if ( USE_REG ) begin : ff_160
        reg   lut_160_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_160_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_160_ff <= lut_160_out;
            end
        end
        
        assign out_data[160] = lut_160_ff;
    end
    else begin : no_ff_160
        assign out_data[160] = lut_160_out;
    end
    endgenerate
    
    
    
    // LUT : 161
    wire [15:0] lut_161_table = 16'b0011001101110011;
    wire [3:0] lut_161_select = {
                             in_data[506],
                             in_data[614],
                             in_data[302],
                             in_data[480]};
    
    wire lut_161_out = lut_161_table[lut_161_select];
    
    generate
    if ( USE_REG ) begin : ff_161
        reg   lut_161_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_161_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_161_ff <= lut_161_out;
            end
        end
        
        assign out_data[161] = lut_161_ff;
    end
    else begin : no_ff_161
        assign out_data[161] = lut_161_out;
    end
    endgenerate
    
    
    
    // LUT : 162
    wire [15:0] lut_162_table = 16'b1100010011011100;
    wire [3:0] lut_162_select = {
                             in_data[167],
                             in_data[477],
                             in_data[23],
                             in_data[202]};
    
    wire lut_162_out = lut_162_table[lut_162_select];
    
    generate
    if ( USE_REG ) begin : ff_162
        reg   lut_162_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_162_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_162_ff <= lut_162_out;
            end
        end
        
        assign out_data[162] = lut_162_ff;
    end
    else begin : no_ff_162
        assign out_data[162] = lut_162_out;
    end
    endgenerate
    
    
    
    // LUT : 163
    wire [15:0] lut_163_table = 16'b1100110011001101;
    wire [3:0] lut_163_select = {
                             in_data[15],
                             in_data[583],
                             in_data[233],
                             in_data[173]};
    
    wire lut_163_out = lut_163_table[lut_163_select];
    
    generate
    if ( USE_REG ) begin : ff_163
        reg   lut_163_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_163_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_163_ff <= lut_163_out;
            end
        end
        
        assign out_data[163] = lut_163_ff;
    end
    else begin : no_ff_163
        assign out_data[163] = lut_163_out;
    end
    endgenerate
    
    
    
    // LUT : 164
    wire [15:0] lut_164_table = 16'b1011001000100010;
    wire [3:0] lut_164_select = {
                             in_data[565],
                             in_data[331],
                             in_data[538],
                             in_data[487]};
    
    wire lut_164_out = lut_164_table[lut_164_select];
    
    generate
    if ( USE_REG ) begin : ff_164
        reg   lut_164_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_164_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_164_ff <= lut_164_out;
            end
        end
        
        assign out_data[164] = lut_164_ff;
    end
    else begin : no_ff_164
        assign out_data[164] = lut_164_out;
    end
    endgenerate
    
    
    
    // LUT : 165
    wire [15:0] lut_165_table = 16'b0000000011111010;
    wire [3:0] lut_165_select = {
                             in_data[511],
                             in_data[269],
                             in_data[153],
                             in_data[309]};
    
    wire lut_165_out = lut_165_table[lut_165_select];
    
    generate
    if ( USE_REG ) begin : ff_165
        reg   lut_165_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_165_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_165_ff <= lut_165_out;
            end
        end
        
        assign out_data[165] = lut_165_ff;
    end
    else begin : no_ff_165
        assign out_data[165] = lut_165_out;
    end
    endgenerate
    
    
    
    // LUT : 166
    wire [15:0] lut_166_table = 16'b0000001100000011;
    wire [3:0] lut_166_select = {
                             in_data[231],
                             in_data[305],
                             in_data[627],
                             in_data[418]};
    
    wire lut_166_out = lut_166_table[lut_166_select];
    
    generate
    if ( USE_REG ) begin : ff_166
        reg   lut_166_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_166_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_166_ff <= lut_166_out;
            end
        end
        
        assign out_data[166] = lut_166_ff;
    end
    else begin : no_ff_166
        assign out_data[166] = lut_166_out;
    end
    endgenerate
    
    
    
    // LUT : 167
    wire [15:0] lut_167_table = 16'b0101010101011101;
    wire [3:0] lut_167_select = {
                             in_data[621],
                             in_data[120],
                             in_data[208],
                             in_data[488]};
    
    wire lut_167_out = lut_167_table[lut_167_select];
    
    generate
    if ( USE_REG ) begin : ff_167
        reg   lut_167_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_167_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_167_ff <= lut_167_out;
            end
        end
        
        assign out_data[167] = lut_167_ff;
    end
    else begin : no_ff_167
        assign out_data[167] = lut_167_out;
    end
    endgenerate
    
    
    
    // LUT : 168
    wire [15:0] lut_168_table = 16'b1100100010101000;
    wire [3:0] lut_168_select = {
                             in_data[526],
                             in_data[369],
                             in_data[266],
                             in_data[587]};
    
    wire lut_168_out = lut_168_table[lut_168_select];
    
    generate
    if ( USE_REG ) begin : ff_168
        reg   lut_168_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_168_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_168_ff <= lut_168_out;
            end
        end
        
        assign out_data[168] = lut_168_ff;
    end
    else begin : no_ff_168
        assign out_data[168] = lut_168_out;
    end
    endgenerate
    
    
    
    // LUT : 169
    wire [15:0] lut_169_table = 16'b1100110011111100;
    wire [3:0] lut_169_select = {
                             in_data[339],
                             in_data[592],
                             in_data[347],
                             in_data[11]};
    
    wire lut_169_out = lut_169_table[lut_169_select];
    
    generate
    if ( USE_REG ) begin : ff_169
        reg   lut_169_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_169_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_169_ff <= lut_169_out;
            end
        end
        
        assign out_data[169] = lut_169_ff;
    end
    else begin : no_ff_169
        assign out_data[169] = lut_169_out;
    end
    endgenerate
    
    
    
    // LUT : 170
    wire [15:0] lut_170_table = 16'b0101010100000000;
    wire [3:0] lut_170_select = {
                             in_data[373],
                             in_data[527],
                             in_data[612],
                             in_data[358]};
    
    wire lut_170_out = lut_170_table[lut_170_select];
    
    generate
    if ( USE_REG ) begin : ff_170
        reg   lut_170_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_170_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_170_ff <= lut_170_out;
            end
        end
        
        assign out_data[170] = lut_170_ff;
    end
    else begin : no_ff_170
        assign out_data[170] = lut_170_out;
    end
    endgenerate
    
    
    
    // LUT : 171
    wire [15:0] lut_171_table = 16'b0100010001000100;
    wire [3:0] lut_171_select = {
                             in_data[412],
                             in_data[409],
                             in_data[364],
                             in_data[334]};
    
    wire lut_171_out = lut_171_table[lut_171_select];
    
    generate
    if ( USE_REG ) begin : ff_171
        reg   lut_171_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_171_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_171_ff <= lut_171_out;
            end
        end
        
        assign out_data[171] = lut_171_ff;
    end
    else begin : no_ff_171
        assign out_data[171] = lut_171_out;
    end
    endgenerate
    
    
    
    // LUT : 172
    wire [15:0] lut_172_table = 16'b0101000011110000;
    wire [3:0] lut_172_select = {
                             in_data[289],
                             in_data[377],
                             in_data[367],
                             in_data[396]};
    
    wire lut_172_out = lut_172_table[lut_172_select];
    
    generate
    if ( USE_REG ) begin : ff_172
        reg   lut_172_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_172_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_172_ff <= lut_172_out;
            end
        end
        
        assign out_data[172] = lut_172_ff;
    end
    else begin : no_ff_172
        assign out_data[172] = lut_172_out;
    end
    endgenerate
    
    
    
    // LUT : 173
    wire [15:0] lut_173_table = 16'b0000101110111011;
    wire [3:0] lut_173_select = {
                             in_data[333],
                             in_data[384],
                             in_data[152],
                             in_data[122]};
    
    wire lut_173_out = lut_173_table[lut_173_select];
    
    generate
    if ( USE_REG ) begin : ff_173
        reg   lut_173_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_173_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_173_ff <= lut_173_out;
            end
        end
        
        assign out_data[173] = lut_173_ff;
    end
    else begin : no_ff_173
        assign out_data[173] = lut_173_out;
    end
    endgenerate
    
    
    
    // LUT : 174
    wire [15:0] lut_174_table = 16'b0101000111110101;
    wire [3:0] lut_174_select = {
                             in_data[474],
                             in_data[363],
                             in_data[178],
                             in_data[271]};
    
    wire lut_174_out = lut_174_table[lut_174_select];
    
    generate
    if ( USE_REG ) begin : ff_174
        reg   lut_174_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_174_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_174_ff <= lut_174_out;
            end
        end
        
        assign out_data[174] = lut_174_ff;
    end
    else begin : no_ff_174
        assign out_data[174] = lut_174_out;
    end
    endgenerate
    
    
    
    // LUT : 175
    wire [15:0] lut_175_table = 16'b1100110011001100;
    wire [3:0] lut_175_select = {
                             in_data[43],
                             in_data[539],
                             in_data[124],
                             in_data[256]};
    
    wire lut_175_out = lut_175_table[lut_175_select];
    
    generate
    if ( USE_REG ) begin : ff_175
        reg   lut_175_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_175_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_175_ff <= lut_175_out;
            end
        end
        
        assign out_data[175] = lut_175_ff;
    end
    else begin : no_ff_175
        assign out_data[175] = lut_175_out;
    end
    endgenerate
    
    
    
    // LUT : 176
    wire [15:0] lut_176_table = 16'b0101010011111111;
    wire [3:0] lut_176_select = {
                             in_data[406],
                             in_data[456],
                             in_data[500],
                             in_data[212]};
    
    wire lut_176_out = lut_176_table[lut_176_select];
    
    generate
    if ( USE_REG ) begin : ff_176
        reg   lut_176_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_176_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_176_ff <= lut_176_out;
            end
        end
        
        assign out_data[176] = lut_176_ff;
    end
    else begin : no_ff_176
        assign out_data[176] = lut_176_out;
    end
    endgenerate
    
    
    
    // LUT : 177
    wire [15:0] lut_177_table = 16'b1100110010001100;
    wire [3:0] lut_177_select = {
                             in_data[17],
                             in_data[606],
                             in_data[485],
                             in_data[215]};
    
    wire lut_177_out = lut_177_table[lut_177_select];
    
    generate
    if ( USE_REG ) begin : ff_177
        reg   lut_177_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_177_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_177_ff <= lut_177_out;
            end
        end
        
        assign out_data[177] = lut_177_ff;
    end
    else begin : no_ff_177
        assign out_data[177] = lut_177_out;
    end
    endgenerate
    
    
    
    // LUT : 178
    wire [15:0] lut_178_table = 16'b0100010001000101;
    wire [3:0] lut_178_select = {
                             in_data[564],
                             in_data[216],
                             in_data[442],
                             in_data[435]};
    
    wire lut_178_out = lut_178_table[lut_178_select];
    
    generate
    if ( USE_REG ) begin : ff_178
        reg   lut_178_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_178_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_178_ff <= lut_178_out;
            end
        end
        
        assign out_data[178] = lut_178_ff;
    end
    else begin : no_ff_178
        assign out_data[178] = lut_178_out;
    end
    endgenerate
    
    
    
    // LUT : 179
    wire [15:0] lut_179_table = 16'b0000001000110011;
    wire [3:0] lut_179_select = {
                             in_data[224],
                             in_data[337],
                             in_data[192],
                             in_data[104]};
    
    wire lut_179_out = lut_179_table[lut_179_select];
    
    generate
    if ( USE_REG ) begin : ff_179
        reg   lut_179_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_179_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_179_ff <= lut_179_out;
            end
        end
        
        assign out_data[179] = lut_179_ff;
    end
    else begin : no_ff_179
        assign out_data[179] = lut_179_out;
    end
    endgenerate
    
    
    
    // LUT : 180
    wire [15:0] lut_180_table = 16'b1010001010110010;
    wire [3:0] lut_180_select = {
                             in_data[326],
                             in_data[19],
                             in_data[113],
                             in_data[531]};
    
    wire lut_180_out = lut_180_table[lut_180_select];
    
    generate
    if ( USE_REG ) begin : ff_180
        reg   lut_180_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_180_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_180_ff <= lut_180_out;
            end
        end
        
        assign out_data[180] = lut_180_ff;
    end
    else begin : no_ff_180
        assign out_data[180] = lut_180_out;
    end
    endgenerate
    
    
    
    // LUT : 181
    wire [15:0] lut_181_table = 16'b0000111101011111;
    wire [3:0] lut_181_select = {
                             in_data[290],
                             in_data[187],
                             in_data[566],
                             in_data[35]};
    
    wire lut_181_out = lut_181_table[lut_181_select];
    
    generate
    if ( USE_REG ) begin : ff_181
        reg   lut_181_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_181_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_181_ff <= lut_181_out;
            end
        end
        
        assign out_data[181] = lut_181_ff;
    end
    else begin : no_ff_181
        assign out_data[181] = lut_181_out;
    end
    endgenerate
    
    
    
    // LUT : 182
    wire [15:0] lut_182_table = 16'b0010001000111011;
    wire [3:0] lut_182_select = {
                             in_data[150],
                             in_data[1],
                             in_data[467],
                             in_data[228]};
    
    wire lut_182_out = lut_182_table[lut_182_select];
    
    generate
    if ( USE_REG ) begin : ff_182
        reg   lut_182_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_182_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_182_ff <= lut_182_out;
            end
        end
        
        assign out_data[182] = lut_182_ff;
    end
    else begin : no_ff_182
        assign out_data[182] = lut_182_out;
    end
    endgenerate
    
    
    
    // LUT : 183
    wire [15:0] lut_183_table = 16'b0001000101110111;
    wire [3:0] lut_183_select = {
                             in_data[112],
                             in_data[295],
                             in_data[537],
                             in_data[462]};
    
    wire lut_183_out = lut_183_table[lut_183_select];
    
    generate
    if ( USE_REG ) begin : ff_183
        reg   lut_183_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_183_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_183_ff <= lut_183_out;
            end
        end
        
        assign out_data[183] = lut_183_ff;
    end
    else begin : no_ff_183
        assign out_data[183] = lut_183_out;
    end
    endgenerate
    
    
    
    // LUT : 184
    wire [15:0] lut_184_table = 16'b1111010111110111;
    wire [3:0] lut_184_select = {
                             in_data[610],
                             in_data[482],
                             in_data[628],
                             in_data[620]};
    
    wire lut_184_out = lut_184_table[lut_184_select];
    
    generate
    if ( USE_REG ) begin : ff_184
        reg   lut_184_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_184_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_184_ff <= lut_184_out;
            end
        end
        
        assign out_data[184] = lut_184_ff;
    end
    else begin : no_ff_184
        assign out_data[184] = lut_184_out;
    end
    endgenerate
    
    
    
    // LUT : 185
    wire [15:0] lut_185_table = 16'b0100010101011111;
    wire [3:0] lut_185_select = {
                             in_data[92],
                             in_data[342],
                             in_data[300],
                             in_data[572]};
    
    wire lut_185_out = lut_185_table[lut_185_select];
    
    generate
    if ( USE_REG ) begin : ff_185
        reg   lut_185_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_185_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_185_ff <= lut_185_out;
            end
        end
        
        assign out_data[185] = lut_185_ff;
    end
    else begin : no_ff_185
        assign out_data[185] = lut_185_out;
    end
    endgenerate
    
    
    
    // LUT : 186
    wire [15:0] lut_186_table = 16'b0111001100010000;
    wire [3:0] lut_186_select = {
                             in_data[204],
                             in_data[542],
                             in_data[574],
                             in_data[524]};
    
    wire lut_186_out = lut_186_table[lut_186_select];
    
    generate
    if ( USE_REG ) begin : ff_186
        reg   lut_186_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_186_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_186_ff <= lut_186_out;
            end
        end
        
        assign out_data[186] = lut_186_ff;
    end
    else begin : no_ff_186
        assign out_data[186] = lut_186_out;
    end
    endgenerate
    
    
    
    // LUT : 187
    wire [15:0] lut_187_table = 16'b0100010011010100;
    wire [3:0] lut_187_select = {
                             in_data[26],
                             in_data[513],
                             in_data[308],
                             in_data[503]};
    
    wire lut_187_out = lut_187_table[lut_187_select];
    
    generate
    if ( USE_REG ) begin : ff_187
        reg   lut_187_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_187_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_187_ff <= lut_187_out;
            end
        end
        
        assign out_data[187] = lut_187_ff;
    end
    else begin : no_ff_187
        assign out_data[187] = lut_187_out;
    end
    endgenerate
    
    
    
    // LUT : 188
    wire [15:0] lut_188_table = 16'b1100110011001100;
    wire [3:0] lut_188_select = {
                             in_data[293],
                             in_data[470],
                             in_data[518],
                             in_data[629]};
    
    wire lut_188_out = lut_188_table[lut_188_select];
    
    generate
    if ( USE_REG ) begin : ff_188
        reg   lut_188_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_188_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_188_ff <= lut_188_out;
            end
        end
        
        assign out_data[188] = lut_188_ff;
    end
    else begin : no_ff_188
        assign out_data[188] = lut_188_out;
    end
    endgenerate
    
    
    
    // LUT : 189
    wire [15:0] lut_189_table = 16'b1011000100110000;
    wire [3:0] lut_189_select = {
                             in_data[21],
                             in_data[444],
                             in_data[516],
                             in_data[283]};
    
    wire lut_189_out = lut_189_table[lut_189_select];
    
    generate
    if ( USE_REG ) begin : ff_189
        reg   lut_189_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_189_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_189_ff <= lut_189_out;
            end
        end
        
        assign out_data[189] = lut_189_ff;
    end
    else begin : no_ff_189
        assign out_data[189] = lut_189_out;
    end
    endgenerate
    
    
    
    // LUT : 190
    wire [15:0] lut_190_table = 16'b0111011111110111;
    wire [3:0] lut_190_select = {
                             in_data[454],
                             in_data[354],
                             in_data[179],
                             in_data[407]};
    
    wire lut_190_out = lut_190_table[lut_190_select];
    
    generate
    if ( USE_REG ) begin : ff_190
        reg   lut_190_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_190_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_190_ff <= lut_190_out;
            end
        end
        
        assign out_data[190] = lut_190_ff;
    end
    else begin : no_ff_190
        assign out_data[190] = lut_190_out;
    end
    endgenerate
    
    
    
    // LUT : 191
    wire [15:0] lut_191_table = 16'b0000000011111111;
    wire [3:0] lut_191_select = {
                             in_data[69],
                             in_data[200],
                             in_data[545],
                             in_data[590]};
    
    wire lut_191_out = lut_191_table[lut_191_select];
    
    generate
    if ( USE_REG ) begin : ff_191
        reg   lut_191_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_191_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_191_ff <= lut_191_out;
            end
        end
        
        assign out_data[191] = lut_191_ff;
    end
    else begin : no_ff_191
        assign out_data[191] = lut_191_out;
    end
    endgenerate
    
    
    
    // LUT : 192
    wire [15:0] lut_192_table = 16'b1100110101001100;
    wire [3:0] lut_192_select = {
                             in_data[162],
                             in_data[429],
                             in_data[630],
                             in_data[54]};
    
    wire lut_192_out = lut_192_table[lut_192_select];
    
    generate
    if ( USE_REG ) begin : ff_192
        reg   lut_192_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_192_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_192_ff <= lut_192_out;
            end
        end
        
        assign out_data[192] = lut_192_ff;
    end
    else begin : no_ff_192
        assign out_data[192] = lut_192_out;
    end
    endgenerate
    
    
    
    // LUT : 193
    wire [15:0] lut_193_table = 16'b1110110010000000;
    wire [3:0] lut_193_select = {
                             in_data[371],
                             in_data[346],
                             in_data[195],
                             in_data[370]};
    
    wire lut_193_out = lut_193_table[lut_193_select];
    
    generate
    if ( USE_REG ) begin : ff_193
        reg   lut_193_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_193_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_193_ff <= lut_193_out;
            end
        end
        
        assign out_data[193] = lut_193_ff;
    end
    else begin : no_ff_193
        assign out_data[193] = lut_193_out;
    end
    endgenerate
    
    
    
    // LUT : 194
    wire [15:0] lut_194_table = 16'b0000010100010101;
    wire [3:0] lut_194_select = {
                             in_data[169],
                             in_data[552],
                             in_data[25],
                             in_data[199]};
    
    wire lut_194_out = lut_194_table[lut_194_select];
    
    generate
    if ( USE_REG ) begin : ff_194
        reg   lut_194_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_194_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_194_ff <= lut_194_out;
            end
        end
        
        assign out_data[194] = lut_194_ff;
    end
    else begin : no_ff_194
        assign out_data[194] = lut_194_out;
    end
    endgenerate
    
    
    
    // LUT : 195
    wire [15:0] lut_195_table = 16'b1101010011111111;
    wire [3:0] lut_195_select = {
                             in_data[413],
                             in_data[157],
                             in_data[495],
                             in_data[555]};
    
    wire lut_195_out = lut_195_table[lut_195_select];
    
    generate
    if ( USE_REG ) begin : ff_195
        reg   lut_195_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_195_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_195_ff <= lut_195_out;
            end
        end
        
        assign out_data[195] = lut_195_ff;
    end
    else begin : no_ff_195
        assign out_data[195] = lut_195_out;
    end
    endgenerate
    
    
    
    // LUT : 196
    wire [15:0] lut_196_table = 16'b1111111100000111;
    wire [3:0] lut_196_select = {
                             in_data[341],
                             in_data[196],
                             in_data[458],
                             in_data[359]};
    
    wire lut_196_out = lut_196_table[lut_196_select];
    
    generate
    if ( USE_REG ) begin : ff_196
        reg   lut_196_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_196_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_196_ff <= lut_196_out;
            end
        end
        
        assign out_data[196] = lut_196_ff;
    end
    else begin : no_ff_196
        assign out_data[196] = lut_196_out;
    end
    endgenerate
    
    
    
    // LUT : 197
    wire [15:0] lut_197_table = 16'b0000010011001110;
    wire [3:0] lut_197_select = {
                             in_data[558],
                             in_data[595],
                             in_data[97],
                             in_data[395]};
    
    wire lut_197_out = lut_197_table[lut_197_select];
    
    generate
    if ( USE_REG ) begin : ff_197
        reg   lut_197_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_197_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_197_ff <= lut_197_out;
            end
        end
        
        assign out_data[197] = lut_197_ff;
    end
    else begin : no_ff_197
        assign out_data[197] = lut_197_out;
    end
    endgenerate
    
    
    
    // LUT : 198
    wire [15:0] lut_198_table = 16'b1111000011110000;
    wire [3:0] lut_198_select = {
                             in_data[240],
                             in_data[291],
                             in_data[568],
                             in_data[533]};
    
    wire lut_198_out = lut_198_table[lut_198_select];
    
    generate
    if ( USE_REG ) begin : ff_198
        reg   lut_198_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_198_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_198_ff <= lut_198_out;
            end
        end
        
        assign out_data[198] = lut_198_ff;
    end
    else begin : no_ff_198
        assign out_data[198] = lut_198_out;
    end
    endgenerate
    
    
    
    // LUT : 199
    wire [15:0] lut_199_table = 16'b1110100011101100;
    wire [3:0] lut_199_select = {
                             in_data[48],
                             in_data[41],
                             in_data[553],
                             in_data[222]};
    
    wire lut_199_out = lut_199_table[lut_199_select];
    
    generate
    if ( USE_REG ) begin : ff_199
        reg   lut_199_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_199_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_199_ff <= lut_199_out;
            end
        end
        
        assign out_data[199] = lut_199_ff;
    end
    else begin : no_ff_199
        assign out_data[199] = lut_199_out;
    end
    endgenerate
    
    
    
    // LUT : 200
    wire [15:0] lut_200_table = 16'b0000001110111111;
    wire [3:0] lut_200_select = {
                             in_data[338],
                             in_data[351],
                             in_data[391],
                             in_data[129]};
    
    wire lut_200_out = lut_200_table[lut_200_select];
    
    generate
    if ( USE_REG ) begin : ff_200
        reg   lut_200_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_200_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_200_ff <= lut_200_out;
            end
        end
        
        assign out_data[200] = lut_200_ff;
    end
    else begin : no_ff_200
        assign out_data[200] = lut_200_out;
    end
    endgenerate
    
    
    
    // LUT : 201
    wire [15:0] lut_201_table = 16'b1100000011000100;
    wire [3:0] lut_201_select = {
                             in_data[519],
                             in_data[479],
                             in_data[306],
                             in_data[138]};
    
    wire lut_201_out = lut_201_table[lut_201_select];
    
    generate
    if ( USE_REG ) begin : ff_201
        reg   lut_201_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_201_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_201_ff <= lut_201_out;
            end
        end
        
        assign out_data[201] = lut_201_ff;
    end
    else begin : no_ff_201
        assign out_data[201] = lut_201_out;
    end
    endgenerate
    
    
    
    // LUT : 202
    wire [15:0] lut_202_table = 16'b0101010100010101;
    wire [3:0] lut_202_select = {
                             in_data[447],
                             in_data[414],
                             in_data[160],
                             in_data[284]};
    
    wire lut_202_out = lut_202_table[lut_202_select];
    
    generate
    if ( USE_REG ) begin : ff_202
        reg   lut_202_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_202_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_202_ff <= lut_202_out;
            end
        end
        
        assign out_data[202] = lut_202_ff;
    end
    else begin : no_ff_202
        assign out_data[202] = lut_202_out;
    end
    endgenerate
    
    
    
    // LUT : 203
    wire [15:0] lut_203_table = 16'b0000010000010011;
    wire [3:0] lut_203_select = {
                             in_data[180],
                             in_data[286],
                             in_data[489],
                             in_data[76]};
    
    wire lut_203_out = lut_203_table[lut_203_select];
    
    generate
    if ( USE_REG ) begin : ff_203
        reg   lut_203_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_203_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_203_ff <= lut_203_out;
            end
        end
        
        assign out_data[203] = lut_203_ff;
    end
    else begin : no_ff_203
        assign out_data[203] = lut_203_out;
    end
    endgenerate
    
    
    
    // LUT : 204
    wire [15:0] lut_204_table = 16'b1010101100100011;
    wire [3:0] lut_204_select = {
                             in_data[64],
                             in_data[163],
                             in_data[410],
                             in_data[101]};
    
    wire lut_204_out = lut_204_table[lut_204_select];
    
    generate
    if ( USE_REG ) begin : ff_204
        reg   lut_204_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_204_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_204_ff <= lut_204_out;
            end
        end
        
        assign out_data[204] = lut_204_ff;
    end
    else begin : no_ff_204
        assign out_data[204] = lut_204_out;
    end
    endgenerate
    
    
    
    // LUT : 205
    wire [15:0] lut_205_table = 16'b0001011100010111;
    wire [3:0] lut_205_select = {
                             in_data[312],
                             in_data[445],
                             in_data[426],
                             in_data[637]};
    
    wire lut_205_out = lut_205_table[lut_205_select];
    
    generate
    if ( USE_REG ) begin : ff_205
        reg   lut_205_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_205_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_205_ff <= lut_205_out;
            end
        end
        
        assign out_data[205] = lut_205_ff;
    end
    else begin : no_ff_205
        assign out_data[205] = lut_205_out;
    end
    endgenerate
    
    
    
    // LUT : 206
    wire [15:0] lut_206_table = 16'b1110110010101000;
    wire [3:0] lut_206_select = {
                             in_data[143],
                             in_data[625],
                             in_data[455],
                             in_data[151]};
    
    wire lut_206_out = lut_206_table[lut_206_select];
    
    generate
    if ( USE_REG ) begin : ff_206
        reg   lut_206_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_206_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_206_ff <= lut_206_out;
            end
        end
        
        assign out_data[206] = lut_206_ff;
    end
    else begin : no_ff_206
        assign out_data[206] = lut_206_out;
    end
    endgenerate
    
    
    
    // LUT : 207
    wire [15:0] lut_207_table = 16'b1100111010001010;
    wire [3:0] lut_207_select = {
                             in_data[144],
                             in_data[175],
                             in_data[415],
                             in_data[299]};
    
    wire lut_207_out = lut_207_table[lut_207_select];
    
    generate
    if ( USE_REG ) begin : ff_207
        reg   lut_207_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_207_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_207_ff <= lut_207_out;
            end
        end
        
        assign out_data[207] = lut_207_ff;
    end
    else begin : no_ff_207
        assign out_data[207] = lut_207_out;
    end
    endgenerate
    
    
    
    // LUT : 208
    wire [15:0] lut_208_table = 16'b1110100011101100;
    wire [3:0] lut_208_select = {
                             in_data[203],
                             in_data[55],
                             in_data[402],
                             in_data[603]};
    
    wire lut_208_out = lut_208_table[lut_208_select];
    
    generate
    if ( USE_REG ) begin : ff_208
        reg   lut_208_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_208_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_208_ff <= lut_208_out;
            end
        end
        
        assign out_data[208] = lut_208_ff;
    end
    else begin : no_ff_208
        assign out_data[208] = lut_208_out;
    end
    endgenerate
    
    
    
    // LUT : 209
    wire [15:0] lut_209_table = 16'b0101111100000101;
    wire [3:0] lut_209_select = {
                             in_data[509],
                             in_data[2],
                             in_data[382],
                             in_data[248]};
    
    wire lut_209_out = lut_209_table[lut_209_select];
    
    generate
    if ( USE_REG ) begin : ff_209
        reg   lut_209_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_209_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_209_ff <= lut_209_out;
            end
        end
        
        assign out_data[209] = lut_209_ff;
    end
    else begin : no_ff_209
        assign out_data[209] = lut_209_out;
    end
    endgenerate
    
    
    
    // LUT : 210
    wire [15:0] lut_210_table = 16'b0000000010001111;
    wire [3:0] lut_210_select = {
                             in_data[322],
                             in_data[438],
                             in_data[83],
                             in_data[514]};
    
    wire lut_210_out = lut_210_table[lut_210_select];
    
    generate
    if ( USE_REG ) begin : ff_210
        reg   lut_210_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_210_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_210_ff <= lut_210_out;
            end
        end
        
        assign out_data[210] = lut_210_ff;
    end
    else begin : no_ff_210
        assign out_data[210] = lut_210_out;
    end
    endgenerate
    
    
    
    // LUT : 211
    wire [15:0] lut_211_table = 16'b0100111101001100;
    wire [3:0] lut_211_select = {
                             in_data[457],
                             in_data[490],
                             in_data[66],
                             in_data[381]};
    
    wire lut_211_out = lut_211_table[lut_211_select];
    
    generate
    if ( USE_REG ) begin : ff_211
        reg   lut_211_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_211_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_211_ff <= lut_211_out;
            end
        end
        
        assign out_data[211] = lut_211_ff;
    end
    else begin : no_ff_211
        assign out_data[211] = lut_211_out;
    end
    endgenerate
    
    
    
    // LUT : 212
    wire [15:0] lut_212_table = 16'b1101110101010100;
    wire [3:0] lut_212_select = {
                             in_data[185],
                             in_data[401],
                             in_data[298],
                             in_data[99]};
    
    wire lut_212_out = lut_212_table[lut_212_select];
    
    generate
    if ( USE_REG ) begin : ff_212
        reg   lut_212_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_212_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_212_ff <= lut_212_out;
            end
        end
        
        assign out_data[212] = lut_212_ff;
    end
    else begin : no_ff_212
        assign out_data[212] = lut_212_out;
    end
    endgenerate
    
    
    
    // LUT : 213
    wire [15:0] lut_213_table = 16'b0000000011111111;
    wire [3:0] lut_213_select = {
                             in_data[237],
                             in_data[265],
                             in_data[98],
                             in_data[523]};
    
    wire lut_213_out = lut_213_table[lut_213_select];
    
    generate
    if ( USE_REG ) begin : ff_213
        reg   lut_213_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_213_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_213_ff <= lut_213_out;
            end
        end
        
        assign out_data[213] = lut_213_ff;
    end
    else begin : no_ff_213
        assign out_data[213] = lut_213_out;
    end
    endgenerate
    
    
    
    // LUT : 214
    wire [15:0] lut_214_table = 16'b1101111101001100;
    wire [3:0] lut_214_select = {
                             in_data[344],
                             in_data[602],
                             in_data[343],
                             in_data[235]};
    
    wire lut_214_out = lut_214_table[lut_214_select];
    
    generate
    if ( USE_REG ) begin : ff_214
        reg   lut_214_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_214_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_214_ff <= lut_214_out;
            end
        end
        
        assign out_data[214] = lut_214_ff;
    end
    else begin : no_ff_214
        assign out_data[214] = lut_214_out;
    end
    endgenerate
    
    
    
    // LUT : 215
    wire [15:0] lut_215_table = 16'b0100110001001111;
    wire [3:0] lut_215_select = {
                             in_data[548],
                             in_data[605],
                             in_data[349],
                             in_data[634]};
    
    wire lut_215_out = lut_215_table[lut_215_select];
    
    generate
    if ( USE_REG ) begin : ff_215
        reg   lut_215_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_215_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_215_ff <= lut_215_out;
            end
        end
        
        assign out_data[215] = lut_215_ff;
    end
    else begin : no_ff_215
        assign out_data[215] = lut_215_out;
    end
    endgenerate
    
    
    
    // LUT : 216
    wire [15:0] lut_216_table = 16'b1111010001000000;
    wire [3:0] lut_216_select = {
                             in_data[465],
                             in_data[130],
                             in_data[255],
                             in_data[89]};
    
    wire lut_216_out = lut_216_table[lut_216_select];
    
    generate
    if ( USE_REG ) begin : ff_216
        reg   lut_216_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_216_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_216_ff <= lut_216_out;
            end
        end
        
        assign out_data[216] = lut_216_ff;
    end
    else begin : no_ff_216
        assign out_data[216] = lut_216_out;
    end
    endgenerate
    
    
    
    // LUT : 217
    wire [15:0] lut_217_table = 16'b1010111110101010;
    wire [3:0] lut_217_select = {
                             in_data[471],
                             in_data[596],
                             in_data[194],
                             in_data[582]};
    
    wire lut_217_out = lut_217_table[lut_217_select];
    
    generate
    if ( USE_REG ) begin : ff_217
        reg   lut_217_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_217_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_217_ff <= lut_217_out;
            end
        end
        
        assign out_data[217] = lut_217_ff;
    end
    else begin : no_ff_217
        assign out_data[217] = lut_217_out;
    end
    endgenerate
    
    
    
    // LUT : 218
    wire [15:0] lut_218_table = 16'b1000010011001100;
    wire [3:0] lut_218_select = {
                             in_data[218],
                             in_data[90],
                             in_data[608],
                             in_data[588]};
    
    wire lut_218_out = lut_218_table[lut_218_select];
    
    generate
    if ( USE_REG ) begin : ff_218
        reg   lut_218_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_218_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_218_ff <= lut_218_out;
            end
        end
        
        assign out_data[218] = lut_218_ff;
    end
    else begin : no_ff_218
        assign out_data[218] = lut_218_out;
    end
    endgenerate
    
    
    
    // LUT : 219
    wire [15:0] lut_219_table = 16'b1110111010000000;
    wire [3:0] lut_219_select = {
                             in_data[374],
                             in_data[546],
                             in_data[205],
                             in_data[51]};
    
    wire lut_219_out = lut_219_table[lut_219_select];
    
    generate
    if ( USE_REG ) begin : ff_219
        reg   lut_219_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_219_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_219_ff <= lut_219_out;
            end
        end
        
        assign out_data[219] = lut_219_ff;
    end
    else begin : no_ff_219
        assign out_data[219] = lut_219_out;
    end
    endgenerate
    
    
    
    // LUT : 220
    wire [15:0] lut_220_table = 16'b0000111111111111;
    wire [3:0] lut_220_select = {
                             in_data[77],
                             in_data[601],
                             in_data[521],
                             in_data[5]};
    
    wire lut_220_out = lut_220_table[lut_220_select];
    
    generate
    if ( USE_REG ) begin : ff_220
        reg   lut_220_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_220_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_220_ff <= lut_220_out;
            end
        end
        
        assign out_data[220] = lut_220_ff;
    end
    else begin : no_ff_220
        assign out_data[220] = lut_220_out;
    end
    endgenerate
    
    
    
    // LUT : 221
    wire [15:0] lut_221_table = 16'b0001011100000101;
    wire [3:0] lut_221_select = {
                             in_data[8],
                             in_data[310],
                             in_data[247],
                             in_data[464]};
    
    wire lut_221_out = lut_221_table[lut_221_select];
    
    generate
    if ( USE_REG ) begin : ff_221
        reg   lut_221_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_221_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_221_ff <= lut_221_out;
            end
        end
        
        assign out_data[221] = lut_221_ff;
    end
    else begin : no_ff_221
        assign out_data[221] = lut_221_out;
    end
    endgenerate
    
    
    
    // LUT : 222
    wire [15:0] lut_222_table = 16'b1100110000000000;
    wire [3:0] lut_222_select = {
                             in_data[615],
                             in_data[221],
                             in_data[109],
                             in_data[183]};
    
    wire lut_222_out = lut_222_table[lut_222_select];
    
    generate
    if ( USE_REG ) begin : ff_222
        reg   lut_222_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_222_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_222_ff <= lut_222_out;
            end
        end
        
        assign out_data[222] = lut_222_ff;
    end
    else begin : no_ff_222
        assign out_data[222] = lut_222_out;
    end
    endgenerate
    
    
    
    // LUT : 223
    wire [15:0] lut_223_table = 16'b1000100010001110;
    wire [3:0] lut_223_select = {
                             in_data[146],
                             in_data[107],
                             in_data[356],
                             in_data[174]};
    
    wire lut_223_out = lut_223_table[lut_223_select];
    
    generate
    if ( USE_REG ) begin : ff_223
        reg   lut_223_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_223_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_223_ff <= lut_223_out;
            end
        end
        
        assign out_data[223] = lut_223_ff;
    end
    else begin : no_ff_223
        assign out_data[223] = lut_223_out;
    end
    endgenerate
    
    
    
    // LUT : 224
    wire [15:0] lut_224_table = 16'b0111011101010100;
    wire [3:0] lut_224_select = {
                             in_data[379],
                             in_data[619],
                             in_data[313],
                             in_data[376]};
    
    wire lut_224_out = lut_224_table[lut_224_select];
    
    generate
    if ( USE_REG ) begin : ff_224
        reg   lut_224_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_224_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_224_ff <= lut_224_out;
            end
        end
        
        assign out_data[224] = lut_224_ff;
    end
    else begin : no_ff_224
        assign out_data[224] = lut_224_out;
    end
    endgenerate
    
    
    
    // LUT : 225
    wire [15:0] lut_225_table = 16'b0010001000110011;
    wire [3:0] lut_225_select = {
                             in_data[188],
                             in_data[473],
                             in_data[557],
                             in_data[281]};
    
    wire lut_225_out = lut_225_table[lut_225_select];
    
    generate
    if ( USE_REG ) begin : ff_225
        reg   lut_225_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_225_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_225_ff <= lut_225_out;
            end
        end
        
        assign out_data[225] = lut_225_ff;
    end
    else begin : no_ff_225
        assign out_data[225] = lut_225_out;
    end
    endgenerate
    
    
    
    // LUT : 226
    wire [15:0] lut_226_table = 16'b1110010011110100;
    wire [3:0] lut_226_select = {
                             in_data[9],
                             in_data[393],
                             in_data[505],
                             in_data[176]};
    
    wire lut_226_out = lut_226_table[lut_226_select];
    
    generate
    if ( USE_REG ) begin : ff_226
        reg   lut_226_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_226_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_226_ff <= lut_226_out;
            end
        end
        
        assign out_data[226] = lut_226_ff;
    end
    else begin : no_ff_226
        assign out_data[226] = lut_226_out;
    end
    endgenerate
    
    
    
    // LUT : 227
    wire [15:0] lut_227_table = 16'b1010000010110010;
    wire [3:0] lut_227_select = {
                             in_data[534],
                             in_data[448],
                             in_data[133],
                             in_data[139]};
    
    wire lut_227_out = lut_227_table[lut_227_select];
    
    generate
    if ( USE_REG ) begin : ff_227
        reg   lut_227_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_227_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_227_ff <= lut_227_out;
            end
        end
        
        assign out_data[227] = lut_227_ff;
    end
    else begin : no_ff_227
        assign out_data[227] = lut_227_out;
    end
    endgenerate
    
    
    
    // LUT : 228
    wire [15:0] lut_228_table = 16'b1011001100110010;
    wire [3:0] lut_228_select = {
                             in_data[361],
                             in_data[206],
                             in_data[626],
                             in_data[241]};
    
    wire lut_228_out = lut_228_table[lut_228_select];
    
    generate
    if ( USE_REG ) begin : ff_228
        reg   lut_228_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_228_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_228_ff <= lut_228_out;
            end
        end
        
        assign out_data[228] = lut_228_ff;
    end
    else begin : no_ff_228
        assign out_data[228] = lut_228_out;
    end
    endgenerate
    
    
    
    // LUT : 229
    wire [15:0] lut_229_table = 16'b0010001010101010;
    wire [3:0] lut_229_select = {
                             in_data[123],
                             in_data[633],
                             in_data[128],
                             in_data[125]};
    
    wire lut_229_out = lut_229_table[lut_229_select];
    
    generate
    if ( USE_REG ) begin : ff_229
        reg   lut_229_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_229_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_229_ff <= lut_229_out;
            end
        end
        
        assign out_data[229] = lut_229_ff;
    end
    else begin : no_ff_229
        assign out_data[229] = lut_229_out;
    end
    endgenerate
    
    
    
    // LUT : 230
    wire [15:0] lut_230_table = 16'b0011001100110111;
    wire [3:0] lut_230_select = {
                             in_data[554],
                             in_data[436],
                             in_data[14],
                             in_data[148]};
    
    wire lut_230_out = lut_230_table[lut_230_select];
    
    generate
    if ( USE_REG ) begin : ff_230
        reg   lut_230_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_230_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_230_ff <= lut_230_out;
            end
        end
        
        assign out_data[230] = lut_230_ff;
    end
    else begin : no_ff_230
        assign out_data[230] = lut_230_out;
    end
    endgenerate
    
    
    
    // LUT : 231
    wire [15:0] lut_231_table = 16'b1111000011110010;
    wire [3:0] lut_231_select = {
                             in_data[400],
                             in_data[451],
                             in_data[589],
                             in_data[323]};
    
    wire lut_231_out = lut_231_table[lut_231_select];
    
    generate
    if ( USE_REG ) begin : ff_231
        reg   lut_231_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_231_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_231_ff <= lut_231_out;
            end
        end
        
        assign out_data[231] = lut_231_ff;
    end
    else begin : no_ff_231
        assign out_data[231] = lut_231_out;
    end
    endgenerate
    
    
    
    // LUT : 232
    wire [15:0] lut_232_table = 16'b0101010101010101;
    wire [3:0] lut_232_select = {
                             in_data[461],
                             in_data[168],
                             in_data[74],
                             in_data[106]};
    
    wire lut_232_out = lut_232_table[lut_232_select];
    
    generate
    if ( USE_REG ) begin : ff_232
        reg   lut_232_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_232_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_232_ff <= lut_232_out;
            end
        end
        
        assign out_data[232] = lut_232_ff;
    end
    else begin : no_ff_232
        assign out_data[232] = lut_232_out;
    end
    endgenerate
    
    
    
    // LUT : 233
    wire [15:0] lut_233_table = 16'b0010100011100000;
    wire [3:0] lut_233_select = {
                             in_data[385],
                             in_data[282],
                             in_data[632],
                             in_data[0]};
    
    wire lut_233_out = lut_233_table[lut_233_select];
    
    generate
    if ( USE_REG ) begin : ff_233
        reg   lut_233_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_233_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_233_ff <= lut_233_out;
            end
        end
        
        assign out_data[233] = lut_233_ff;
    end
    else begin : no_ff_233
        assign out_data[233] = lut_233_out;
    end
    endgenerate
    
    
    
    // LUT : 234
    wire [15:0] lut_234_table = 16'b0000000011110000;
    wire [3:0] lut_234_select = {
                             in_data[262],
                             in_data[257],
                             in_data[280],
                             in_data[186]};
    
    wire lut_234_out = lut_234_table[lut_234_select];
    
    generate
    if ( USE_REG ) begin : ff_234
        reg   lut_234_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_234_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_234_ff <= lut_234_out;
            end
        end
        
        assign out_data[234] = lut_234_ff;
    end
    else begin : no_ff_234
        assign out_data[234] = lut_234_out;
    end
    endgenerate
    
    
    
    // LUT : 235
    wire [15:0] lut_235_table = 16'b0000001000101010;
    wire [3:0] lut_235_select = {
                             in_data[198],
                             in_data[631],
                             in_data[484],
                             in_data[131]};
    
    wire lut_235_out = lut_235_table[lut_235_select];
    
    generate
    if ( USE_REG ) begin : ff_235
        reg   lut_235_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_235_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_235_ff <= lut_235_out;
            end
        end
        
        assign out_data[235] = lut_235_ff;
    end
    else begin : no_ff_235
        assign out_data[235] = lut_235_out;
    end
    endgenerate
    
    
    
    // LUT : 236
    wire [15:0] lut_236_table = 16'b1000111010001110;
    wire [3:0] lut_236_select = {
                             in_data[60],
                             in_data[498],
                             in_data[304],
                             in_data[551]};
    
    wire lut_236_out = lut_236_table[lut_236_select];
    
    generate
    if ( USE_REG ) begin : ff_236
        reg   lut_236_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_236_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_236_ff <= lut_236_out;
            end
        end
        
        assign out_data[236] = lut_236_ff;
    end
    else begin : no_ff_236
        assign out_data[236] = lut_236_out;
    end
    endgenerate
    
    
    
    // LUT : 237
    wire [15:0] lut_237_table = 16'b0100111100000101;
    wire [3:0] lut_237_select = {
                             in_data[108],
                             in_data[159],
                             in_data[12],
                             in_data[201]};
    
    wire lut_237_out = lut_237_table[lut_237_select];
    
    generate
    if ( USE_REG ) begin : ff_237
        reg   lut_237_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_237_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_237_ff <= lut_237_out;
            end
        end
        
        assign out_data[237] = lut_237_ff;
    end
    else begin : no_ff_237
        assign out_data[237] = lut_237_out;
    end
    endgenerate
    
    
    
    // LUT : 238
    wire [15:0] lut_238_table = 16'b1100111100000100;
    wire [3:0] lut_238_select = {
                             in_data[317],
                             in_data[18],
                             in_data[556],
                             in_data[115]};
    
    wire lut_238_out = lut_238_table[lut_238_select];
    
    generate
    if ( USE_REG ) begin : ff_238
        reg   lut_238_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_238_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_238_ff <= lut_238_out;
            end
        end
        
        assign out_data[238] = lut_238_ff;
    end
    else begin : no_ff_238
        assign out_data[238] = lut_238_out;
    end
    endgenerate
    
    
    
    // LUT : 239
    wire [15:0] lut_239_table = 16'b0000001000110011;
    wire [3:0] lut_239_select = {
                             in_data[145],
                             in_data[586],
                             in_data[604],
                             in_data[316]};
    
    wire lut_239_out = lut_239_table[lut_239_select];
    
    generate
    if ( USE_REG ) begin : ff_239
        reg   lut_239_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_239_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_239_ff <= lut_239_out;
            end
        end
        
        assign out_data[239] = lut_239_ff;
    end
    else begin : no_ff_239
        assign out_data[239] = lut_239_out;
    end
    endgenerate
    
    
    
    // LUT : 240
    wire [15:0] lut_240_table = 16'b1010101110101010;
    wire [3:0] lut_240_select = {
                             in_data[86],
                             in_data[190],
                             in_data[261],
                             in_data[184]};
    
    wire lut_240_out = lut_240_table[lut_240_select];
    
    generate
    if ( USE_REG ) begin : ff_240
        reg   lut_240_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_240_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_240_ff <= lut_240_out;
            end
        end
        
        assign out_data[240] = lut_240_ff;
    end
    else begin : no_ff_240
        assign out_data[240] = lut_240_out;
    end
    endgenerate
    
    
    
    // LUT : 241
    wire [15:0] lut_241_table = 16'b0000000001010001;
    wire [3:0] lut_241_select = {
                             in_data[57],
                             in_data[264],
                             in_data[353],
                             in_data[622]};
    
    wire lut_241_out = lut_241_table[lut_241_select];
    
    generate
    if ( USE_REG ) begin : ff_241
        reg   lut_241_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_241_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_241_ff <= lut_241_out;
            end
        end
        
        assign out_data[241] = lut_241_ff;
    end
    else begin : no_ff_241
        assign out_data[241] = lut_241_out;
    end
    endgenerate
    
    
    
    // LUT : 242
    wire [15:0] lut_242_table = 16'b0111111100001111;
    wire [3:0] lut_242_select = {
                             in_data[31],
                             in_data[4],
                             in_data[37],
                             in_data[177]};
    
    wire lut_242_out = lut_242_table[lut_242_select];
    
    generate
    if ( USE_REG ) begin : ff_242
        reg   lut_242_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_242_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_242_ff <= lut_242_out;
            end
        end
        
        assign out_data[242] = lut_242_ff;
    end
    else begin : no_ff_242
        assign out_data[242] = lut_242_out;
    end
    endgenerate
    
    
    
    // LUT : 243
    wire [15:0] lut_243_table = 16'b0010101110101111;
    wire [3:0] lut_243_select = {
                             in_data[549],
                             in_data[397],
                             in_data[268],
                             in_data[242]};
    
    wire lut_243_out = lut_243_table[lut_243_select];
    
    generate
    if ( USE_REG ) begin : ff_243
        reg   lut_243_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_243_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_243_ff <= lut_243_out;
            end
        end
        
        assign out_data[243] = lut_243_ff;
    end
    else begin : no_ff_243
        assign out_data[243] = lut_243_out;
    end
    endgenerate
    
    
    
    // LUT : 244
    wire [15:0] lut_244_table = 16'b0000111110111111;
    wire [3:0] lut_244_select = {
                             in_data[501],
                             in_data[78],
                             in_data[253],
                             in_data[81]};
    
    wire lut_244_out = lut_244_table[lut_244_select];
    
    generate
    if ( USE_REG ) begin : ff_244
        reg   lut_244_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_244_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_244_ff <= lut_244_out;
            end
        end
        
        assign out_data[244] = lut_244_ff;
    end
    else begin : no_ff_244
        assign out_data[244] = lut_244_out;
    end
    endgenerate
    
    
    
    // LUT : 245
    wire [15:0] lut_245_table = 16'b0101111100000100;
    wire [3:0] lut_245_select = {
                             in_data[100],
                             in_data[191],
                             in_data[217],
                             in_data[386]};
    
    wire lut_245_out = lut_245_table[lut_245_select];
    
    generate
    if ( USE_REG ) begin : ff_245
        reg   lut_245_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_245_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_245_ff <= lut_245_out;
            end
        end
        
        assign out_data[245] = lut_245_ff;
    end
    else begin : no_ff_245
        assign out_data[245] = lut_245_out;
    end
    endgenerate
    
    
    
    // LUT : 246
    wire [15:0] lut_246_table = 16'b0100111100000101;
    wire [3:0] lut_246_select = {
                             in_data[529],
                             in_data[102],
                             in_data[504],
                             in_data[563]};
    
    wire lut_246_out = lut_246_table[lut_246_select];
    
    generate
    if ( USE_REG ) begin : ff_246
        reg   lut_246_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_246_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_246_ff <= lut_246_out;
            end
        end
        
        assign out_data[246] = lut_246_ff;
    end
    else begin : no_ff_246
        assign out_data[246] = lut_246_out;
    end
    endgenerate
    
    
    
    // LUT : 247
    wire [15:0] lut_247_table = 16'b1101111100001111;
    wire [3:0] lut_247_select = {
                             in_data[497],
                             in_data[278],
                             in_data[91],
                             in_data[223]};
    
    wire lut_247_out = lut_247_table[lut_247_select];
    
    generate
    if ( USE_REG ) begin : ff_247
        reg   lut_247_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_247_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_247_ff <= lut_247_out;
            end
        end
        
        assign out_data[247] = lut_247_ff;
    end
    else begin : no_ff_247
        assign out_data[247] = lut_247_out;
    end
    endgenerate
    
    
    
    // LUT : 248
    wire [15:0] lut_248_table = 16'b1101110011011101;
    wire [3:0] lut_248_select = {
                             in_data[434],
                             in_data[33],
                             in_data[611],
                             in_data[46]};
    
    wire lut_248_out = lut_248_table[lut_248_select];
    
    generate
    if ( USE_REG ) begin : ff_248
        reg   lut_248_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_248_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_248_ff <= lut_248_out;
            end
        end
        
        assign out_data[248] = lut_248_ff;
    end
    else begin : no_ff_248
        assign out_data[248] = lut_248_out;
    end
    endgenerate
    
    
    
    // LUT : 249
    wire [15:0] lut_249_table = 16'b1101010011110100;
    wire [3:0] lut_249_select = {
                             in_data[535],
                             in_data[577],
                             in_data[493],
                             in_data[126]};
    
    wire lut_249_out = lut_249_table[lut_249_select];
    
    generate
    if ( USE_REG ) begin : ff_249
        reg   lut_249_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_249_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_249_ff <= lut_249_out;
            end
        end
        
        assign out_data[249] = lut_249_ff;
    end
    else begin : no_ff_249
        assign out_data[249] = lut_249_out;
    end
    endgenerate
    
    
    
    // LUT : 250
    wire [15:0] lut_250_table = 16'b1100111011001111;
    wire [3:0] lut_250_select = {
                             in_data[491],
                             in_data[79],
                             in_data[36],
                             in_data[460]};
    
    wire lut_250_out = lut_250_table[lut_250_select];
    
    generate
    if ( USE_REG ) begin : ff_250
        reg   lut_250_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_250_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_250_ff <= lut_250_out;
            end
        end
        
        assign out_data[250] = lut_250_ff;
    end
    else begin : no_ff_250
        assign out_data[250] = lut_250_out;
    end
    endgenerate
    
    
    
    // LUT : 251
    wire [15:0] lut_251_table = 16'b1110010011101111;
    wire [3:0] lut_251_select = {
                             in_data[547],
                             in_data[450],
                             in_data[517],
                             in_data[210]};
    
    wire lut_251_out = lut_251_table[lut_251_select];
    
    generate
    if ( USE_REG ) begin : ff_251
        reg   lut_251_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_251_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_251_ff <= lut_251_out;
            end
        end
        
        assign out_data[251] = lut_251_ff;
    end
    else begin : no_ff_251
        assign out_data[251] = lut_251_out;
    end
    endgenerate
    
    
    
    // LUT : 252
    wire [15:0] lut_252_table = 16'b0101010101010101;
    wire [3:0] lut_252_select = {
                             in_data[387],
                             in_data[49],
                             in_data[431],
                             in_data[638]};
    
    wire lut_252_out = lut_252_table[lut_252_select];
    
    generate
    if ( USE_REG ) begin : ff_252
        reg   lut_252_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_252_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_252_ff <= lut_252_out;
            end
        end
        
        assign out_data[252] = lut_252_ff;
    end
    else begin : no_ff_252
        assign out_data[252] = lut_252_out;
    end
    endgenerate
    
    
    
    // LUT : 253
    wire [15:0] lut_253_table = 16'b1000110011001110;
    wire [3:0] lut_253_select = {
                             in_data[425],
                             in_data[368],
                             in_data[296],
                             in_data[567]};
    
    wire lut_253_out = lut_253_table[lut_253_select];
    
    generate
    if ( USE_REG ) begin : ff_253
        reg   lut_253_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_253_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_253_ff <= lut_253_out;
            end
        end
        
        assign out_data[253] = lut_253_ff;
    end
    else begin : no_ff_253
        assign out_data[253] = lut_253_out;
    end
    endgenerate
    
    
    
    // LUT : 254
    wire [15:0] lut_254_table = 16'b0001011100010111;
    wire [3:0] lut_254_select = {
                             in_data[439],
                             in_data[238],
                             in_data[29],
                             in_data[392]};
    
    wire lut_254_out = lut_254_table[lut_254_select];
    
    generate
    if ( USE_REG ) begin : ff_254
        reg   lut_254_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_254_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_254_ff <= lut_254_out;
            end
        end
        
        assign out_data[254] = lut_254_ff;
    end
    else begin : no_ff_254
        assign out_data[254] = lut_254_out;
    end
    endgenerate
    
    
    
    // LUT : 255
    wire [15:0] lut_255_table = 16'b1100000011000000;
    wire [3:0] lut_255_select = {
                             in_data[475],
                             in_data[335],
                             in_data[559],
                             in_data[249]};
    
    wire lut_255_out = lut_255_table[lut_255_select];
    
    generate
    if ( USE_REG ) begin : ff_255
        reg   lut_255_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_255_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_255_ff <= lut_255_out;
            end
        end
        
        assign out_data[255] = lut_255_ff;
    end
    else begin : no_ff_255
        assign out_data[255] = lut_255_out;
    end
    endgenerate
    
    
    
    // LUT : 256
    wire [15:0] lut_256_table = 16'b0000110011001101;
    wire [3:0] lut_256_select = {
                             in_data[576],
                             in_data[52],
                             in_data[544],
                             in_data[61]};
    
    wire lut_256_out = lut_256_table[lut_256_select];
    
    generate
    if ( USE_REG ) begin : ff_256
        reg   lut_256_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_256_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_256_ff <= lut_256_out;
            end
        end
        
        assign out_data[256] = lut_256_ff;
    end
    else begin : no_ff_256
        assign out_data[256] = lut_256_out;
    end
    endgenerate
    
    
    
    // LUT : 257
    wire [15:0] lut_257_table = 16'b1111111100001111;
    wire [3:0] lut_257_select = {
                             in_data[319],
                             in_data[117],
                             in_data[16],
                             in_data[272]};
    
    wire lut_257_out = lut_257_table[lut_257_select];
    
    generate
    if ( USE_REG ) begin : ff_257
        reg   lut_257_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_257_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_257_ff <= lut_257_out;
            end
        end
        
        assign out_data[257] = lut_257_ff;
    end
    else begin : no_ff_257
        assign out_data[257] = lut_257_out;
    end
    endgenerate
    
    
    
    // LUT : 258
    wire [15:0] lut_258_table = 16'b0000110010001110;
    wire [3:0] lut_258_select = {
                             in_data[70],
                             in_data[225],
                             in_data[32],
                             in_data[609]};
    
    wire lut_258_out = lut_258_table[lut_258_select];
    
    generate
    if ( USE_REG ) begin : ff_258
        reg   lut_258_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_258_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_258_ff <= lut_258_out;
            end
        end
        
        assign out_data[258] = lut_258_ff;
    end
    else begin : no_ff_258
        assign out_data[258] = lut_258_out;
    end
    endgenerate
    
    
    
    // LUT : 259
    wire [15:0] lut_259_table = 16'b0010001100110011;
    wire [3:0] lut_259_select = {
                             in_data[562],
                             in_data[580],
                             in_data[383],
                             in_data[42]};
    
    wire lut_259_out = lut_259_table[lut_259_select];
    
    generate
    if ( USE_REG ) begin : ff_259
        reg   lut_259_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_259_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_259_ff <= lut_259_out;
            end
        end
        
        assign out_data[259] = lut_259_ff;
    end
    else begin : no_ff_259
        assign out_data[259] = lut_259_out;
    end
    endgenerate
    
    
    
    // LUT : 260
    wire [15:0] lut_260_table = 16'b1111110011000000;
    wire [3:0] lut_260_select = {
                             in_data[95],
                             in_data[593],
                             in_data[259],
                             in_data[616]};
    
    wire lut_260_out = lut_260_table[lut_260_select];
    
    generate
    if ( USE_REG ) begin : ff_260
        reg   lut_260_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_260_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_260_ff <= lut_260_out;
            end
        end
        
        assign out_data[260] = lut_260_ff;
    end
    else begin : no_ff_260
        assign out_data[260] = lut_260_out;
    end
    endgenerate
    
    
    
    // LUT : 261
    wire [15:0] lut_261_table = 16'b1010101010001010;
    wire [3:0] lut_261_select = {
                             in_data[75],
                             in_data[147],
                             in_data[449],
                             in_data[599]};
    
    wire lut_261_out = lut_261_table[lut_261_select];
    
    generate
    if ( USE_REG ) begin : ff_261
        reg   lut_261_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_261_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_261_ff <= lut_261_out;
            end
        end
        
        assign out_data[261] = lut_261_ff;
    end
    else begin : no_ff_261
        assign out_data[261] = lut_261_out;
    end
    endgenerate
    
    
    
    // LUT : 262
    wire [15:0] lut_262_table = 16'b1010111100001000;
    wire [3:0] lut_262_select = {
                             in_data[244],
                             in_data[229],
                             in_data[132],
                             in_data[294]};
    
    wire lut_262_out = lut_262_table[lut_262_select];
    
    generate
    if ( USE_REG ) begin : ff_262
        reg   lut_262_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_262_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_262_ff <= lut_262_out;
            end
        end
        
        assign out_data[262] = lut_262_ff;
    end
    else begin : no_ff_262
        assign out_data[262] = lut_262_out;
    end
    endgenerate
    
    
    
    // LUT : 263
    wire [15:0] lut_263_table = 16'b1100110011111111;
    wire [3:0] lut_263_select = {
                             in_data[348],
                             in_data[598],
                             in_data[230],
                             in_data[571]};
    
    wire lut_263_out = lut_263_table[lut_263_select];
    
    generate
    if ( USE_REG ) begin : ff_263
        reg   lut_263_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_263_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_263_ff <= lut_263_out;
            end
        end
        
        assign out_data[263] = lut_263_ff;
    end
    else begin : no_ff_263
        assign out_data[263] = lut_263_out;
    end
    endgenerate
    
    
    
    // LUT : 264
    wire [15:0] lut_264_table = 16'b1111110011101000;
    wire [3:0] lut_264_select = {
                             in_data[7],
                             in_data[543],
                             in_data[419],
                             in_data[466]};
    
    wire lut_264_out = lut_264_table[lut_264_select];
    
    generate
    if ( USE_REG ) begin : ff_264
        reg   lut_264_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_264_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_264_ff <= lut_264_out;
            end
        end
        
        assign out_data[264] = lut_264_ff;
    end
    else begin : no_ff_264
        assign out_data[264] = lut_264_out;
    end
    endgenerate
    
    
    
    // LUT : 265
    wire [15:0] lut_265_table = 16'b1100010011000000;
    wire [3:0] lut_265_select = {
                             in_data[440],
                             in_data[352],
                             in_data[22],
                             in_data[20]};
    
    wire lut_265_out = lut_265_table[lut_265_select];
    
    generate
    if ( USE_REG ) begin : ff_265
        reg   lut_265_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_265_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_265_ff <= lut_265_out;
            end
        end
        
        assign out_data[265] = lut_265_ff;
    end
    else begin : no_ff_265
        assign out_data[265] = lut_265_out;
    end
    endgenerate
    
    
    
    // LUT : 266
    wire [15:0] lut_266_table = 16'b1111110011111100;
    wire [3:0] lut_266_select = {
                             in_data[260],
                             in_data[245],
                             in_data[607],
                             in_data[428]};
    
    wire lut_266_out = lut_266_table[lut_266_select];
    
    generate
    if ( USE_REG ) begin : ff_266
        reg   lut_266_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_266_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_266_ff <= lut_266_out;
            end
        end
        
        assign out_data[266] = lut_266_ff;
    end
    else begin : no_ff_266
        assign out_data[266] = lut_266_out;
    end
    endgenerate
    
    
    
    // LUT : 267
    wire [15:0] lut_267_table = 16'b0011101110111011;
    wire [3:0] lut_267_select = {
                             in_data[236],
                             in_data[578],
                             in_data[137],
                             in_data[416]};
    
    wire lut_267_out = lut_267_table[lut_267_select];
    
    generate
    if ( USE_REG ) begin : ff_267
        reg   lut_267_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_267_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_267_ff <= lut_267_out;
            end
        end
        
        assign out_data[267] = lut_267_ff;
    end
    else begin : no_ff_267
        assign out_data[267] = lut_267_out;
    end
    endgenerate
    
    
    
    // LUT : 268
    wire [15:0] lut_268_table = 16'b1111111111110000;
    wire [3:0] lut_268_select = {
                             in_data[591],
                             in_data[581],
                             in_data[618],
                             in_data[82]};
    
    wire lut_268_out = lut_268_table[lut_268_select];
    
    generate
    if ( USE_REG ) begin : ff_268
        reg   lut_268_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_268_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_268_ff <= lut_268_out;
            end
        end
        
        assign out_data[268] = lut_268_ff;
    end
    else begin : no_ff_268
        assign out_data[268] = lut_268_out;
    end
    endgenerate
    
    
    
    // LUT : 269
    wire [15:0] lut_269_table = 16'b0011001101111111;
    wire [3:0] lut_269_select = {
                             in_data[536],
                             in_data[88],
                             in_data[105],
                             in_data[579]};
    
    wire lut_269_out = lut_269_table[lut_269_select];
    
    generate
    if ( USE_REG ) begin : ff_269
        reg   lut_269_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_269_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_269_ff <= lut_269_out;
            end
        end
        
        assign out_data[269] = lut_269_ff;
    end
    else begin : no_ff_269
        assign out_data[269] = lut_269_out;
    end
    endgenerate
    
    
    
    // LUT : 270
    wire [15:0] lut_270_table = 16'b0101010111111111;
    wire [3:0] lut_270_select = {
                             in_data[408],
                             in_data[127],
                             in_data[452],
                             in_data[389]};
    
    wire lut_270_out = lut_270_table[lut_270_select];
    
    generate
    if ( USE_REG ) begin : ff_270
        reg   lut_270_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_270_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_270_ff <= lut_270_out;
            end
        end
        
        assign out_data[270] = lut_270_ff;
    end
    else begin : no_ff_270
        assign out_data[270] = lut_270_out;
    end
    endgenerate
    
    
    
    // LUT : 271
    wire [15:0] lut_271_table = 16'b1110101010101010;
    wire [3:0] lut_271_select = {
                             in_data[314],
                             in_data[424],
                             in_data[510],
                             in_data[525]};
    
    wire lut_271_out = lut_271_table[lut_271_select];
    
    generate
    if ( USE_REG ) begin : ff_271
        reg   lut_271_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_271_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_271_ff <= lut_271_out;
            end
        end
        
        assign out_data[271] = lut_271_ff;
    end
    else begin : no_ff_271
        assign out_data[271] = lut_271_out;
    end
    endgenerate
    
    
    
    // LUT : 272
    wire [15:0] lut_272_table = 16'b1010111000001010;
    wire [3:0] lut_272_select = {
                             in_data[315],
                             in_data[404],
                             in_data[24],
                             in_data[372]};
    
    wire lut_272_out = lut_272_table[lut_272_select];
    
    generate
    if ( USE_REG ) begin : ff_272
        reg   lut_272_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_272_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_272_ff <= lut_272_out;
            end
        end
        
        assign out_data[272] = lut_272_ff;
    end
    else begin : no_ff_272
        assign out_data[272] = lut_272_out;
    end
    endgenerate
    
    
    
    // LUT : 273
    wire [15:0] lut_273_table = 16'b0101010101010101;
    wire [3:0] lut_273_select = {
                             in_data[350],
                             in_data[327],
                             in_data[446],
                             in_data[10]};
    
    wire lut_273_out = lut_273_table[lut_273_select];
    
    generate
    if ( USE_REG ) begin : ff_273
        reg   lut_273_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_273_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_273_ff <= lut_273_out;
            end
        end
        
        assign out_data[273] = lut_273_ff;
    end
    else begin : no_ff_273
        assign out_data[273] = lut_273_out;
    end
    endgenerate
    
    
    
    // LUT : 274
    wire [15:0] lut_274_table = 16'b0101000101010001;
    wire [3:0] lut_274_select = {
                             in_data[30],
                             in_data[623],
                             in_data[85],
                             in_data[496]};
    
    wire lut_274_out = lut_274_table[lut_274_select];
    
    generate
    if ( USE_REG ) begin : ff_274
        reg   lut_274_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_274_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_274_ff <= lut_274_out;
            end
        end
        
        assign out_data[274] = lut_274_ff;
    end
    else begin : no_ff_274
        assign out_data[274] = lut_274_out;
    end
    endgenerate
    
    
    
    // LUT : 275
    wire [15:0] lut_275_table = 16'b0101000011110100;
    wire [3:0] lut_275_select = {
                             in_data[380],
                             in_data[332],
                             in_data[492],
                             in_data[297]};
    
    wire lut_275_out = lut_275_table[lut_275_select];
    
    generate
    if ( USE_REG ) begin : ff_275
        reg   lut_275_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_275_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_275_ff <= lut_275_out;
            end
        end
        
        assign out_data[275] = lut_275_ff;
    end
    else begin : no_ff_275
        assign out_data[275] = lut_275_out;
    end
    endgenerate
    
    
    
    // LUT : 276
    wire [15:0] lut_276_table = 16'b1110100011111000;
    wire [3:0] lut_276_select = {
                             in_data[254],
                             in_data[246],
                             in_data[63],
                             in_data[617]};
    
    wire lut_276_out = lut_276_table[lut_276_select];
    
    generate
    if ( USE_REG ) begin : ff_276
        reg   lut_276_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_276_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_276_ff <= lut_276_out;
            end
        end
        
        assign out_data[276] = lut_276_ff;
    end
    else begin : no_ff_276
        assign out_data[276] = lut_276_out;
    end
    endgenerate
    
    
    
    // LUT : 277
    wire [15:0] lut_277_table = 16'b1111000101110000;
    wire [3:0] lut_277_select = {
                             in_data[39],
                             in_data[324],
                             in_data[53],
                             in_data[94]};
    
    wire lut_277_out = lut_277_table[lut_277_select];
    
    generate
    if ( USE_REG ) begin : ff_277
        reg   lut_277_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_277_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_277_ff <= lut_277_out;
            end
        end
        
        assign out_data[277] = lut_277_ff;
    end
    else begin : no_ff_277
        assign out_data[277] = lut_277_out;
    end
    endgenerate
    
    
    
    // LUT : 278
    wire [15:0] lut_278_table = 16'b0000000111111111;
    wire [3:0] lut_278_select = {
                             in_data[430],
                             in_data[219],
                             in_data[378],
                             in_data[243]};
    
    wire lut_278_out = lut_278_table[lut_278_select];
    
    generate
    if ( USE_REG ) begin : ff_278
        reg   lut_278_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_278_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_278_ff <= lut_278_out;
            end
        end
        
        assign out_data[278] = lut_278_ff;
    end
    else begin : no_ff_278
        assign out_data[278] = lut_278_out;
    end
    endgenerate
    
    
    
    // LUT : 279
    wire [15:0] lut_279_table = 16'b1111110011111010;
    wire [3:0] lut_279_select = {
                             in_data[357],
                             in_data[321],
                             in_data[267],
                             in_data[522]};
    
    wire lut_279_out = lut_279_table[lut_279_select];
    
    generate
    if ( USE_REG ) begin : ff_279
        reg   lut_279_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_279_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_279_ff <= lut_279_out;
            end
        end
        
        assign out_data[279] = lut_279_ff;
    end
    else begin : no_ff_279
        assign out_data[279] = lut_279_out;
    end
    endgenerate
    
    
    
    // LUT : 280
    wire [15:0] lut_280_table = 16'b0011111100111111;
    wire [3:0] lut_280_select = {
                             in_data[181],
                             in_data[156],
                             in_data[486],
                             in_data[398]};
    
    wire lut_280_out = lut_280_table[lut_280_select];
    
    generate
    if ( USE_REG ) begin : ff_280
        reg   lut_280_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_280_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_280_ff <= lut_280_out;
            end
        end
        
        assign out_data[280] = lut_280_ff;
    end
    else begin : no_ff_280
        assign out_data[280] = lut_280_out;
    end
    endgenerate
    
    
    
    // LUT : 281
    wire [15:0] lut_281_table = 16'b1000111000001100;
    wire [3:0] lut_281_select = {
                             in_data[158],
                             in_data[481],
                             in_data[80],
                             in_data[44]};
    
    wire lut_281_out = lut_281_table[lut_281_select];
    
    generate
    if ( USE_REG ) begin : ff_281
        reg   lut_281_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_281_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_281_ff <= lut_281_out;
            end
        end
        
        assign out_data[281] = lut_281_ff;
    end
    else begin : no_ff_281
        assign out_data[281] = lut_281_out;
    end
    endgenerate
    
    
    
    // LUT : 282
    wire [15:0] lut_282_table = 16'b0000000011011100;
    wire [3:0] lut_282_select = {
                             in_data[67],
                             in_data[232],
                             in_data[171],
                             in_data[189]};
    
    wire lut_282_out = lut_282_table[lut_282_select];
    
    generate
    if ( USE_REG ) begin : ff_282
        reg   lut_282_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_282_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_282_ff <= lut_282_out;
            end
        end
        
        assign out_data[282] = lut_282_ff;
    end
    else begin : no_ff_282
        assign out_data[282] = lut_282_out;
    end
    endgenerate
    
    
    
    // LUT : 283
    wire [15:0] lut_283_table = 16'b0000111100001111;
    wire [3:0] lut_283_select = {
                             in_data[561],
                             in_data[530],
                             in_data[441],
                             in_data[275]};
    
    wire lut_283_out = lut_283_table[lut_283_select];
    
    generate
    if ( USE_REG ) begin : ff_283
        reg   lut_283_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_283_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_283_ff <= lut_283_out;
            end
        end
        
        assign out_data[283] = lut_283_ff;
    end
    else begin : no_ff_283
        assign out_data[283] = lut_283_out;
    end
    endgenerate
    
    
    
    // LUT : 284
    wire [15:0] lut_284_table = 16'b0000001110111111;
    wire [3:0] lut_284_select = {
                             in_data[65],
                             in_data[427],
                             in_data[585],
                             in_data[355]};
    
    wire lut_284_out = lut_284_table[lut_284_select];
    
    generate
    if ( USE_REG ) begin : ff_284
        reg   lut_284_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_284_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_284_ff <= lut_284_out;
            end
        end
        
        assign out_data[284] = lut_284_ff;
    end
    else begin : no_ff_284
        assign out_data[284] = lut_284_out;
    end
    endgenerate
    
    
    
    // LUT : 285
    wire [15:0] lut_285_table = 16'b1101110101000100;
    wire [3:0] lut_285_select = {
                             in_data[512],
                             in_data[165],
                             in_data[140],
                             in_data[6]};
    
    wire lut_285_out = lut_285_table[lut_285_select];
    
    generate
    if ( USE_REG ) begin : ff_285
        reg   lut_285_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_285_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_285_ff <= lut_285_out;
            end
        end
        
        assign out_data[285] = lut_285_ff;
    end
    else begin : no_ff_285
        assign out_data[285] = lut_285_out;
    end
    endgenerate
    
    
    
    // LUT : 286
    wire [15:0] lut_286_table = 16'b0000101010101110;
    wire [3:0] lut_286_select = {
                             in_data[258],
                             in_data[154],
                             in_data[285],
                             in_data[111]};
    
    wire lut_286_out = lut_286_table[lut_286_select];
    
    generate
    if ( USE_REG ) begin : ff_286
        reg   lut_286_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_286_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_286_ff <= lut_286_out;
            end
        end
        
        assign out_data[286] = lut_286_ff;
    end
    else begin : no_ff_286
        assign out_data[286] = lut_286_out;
    end
    endgenerate
    
    
    
    // LUT : 287
    wire [15:0] lut_287_table = 16'b0011001100110011;
    wire [3:0] lut_287_select = {
                             in_data[520],
                             in_data[72],
                             in_data[155],
                             in_data[320]};
    
    wire lut_287_out = lut_287_table[lut_287_select];
    
    generate
    if ( USE_REG ) begin : ff_287
        reg   lut_287_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_287_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_287_ff <= lut_287_out;
            end
        end
        
        assign out_data[287] = lut_287_ff;
    end
    else begin : no_ff_287
        assign out_data[287] = lut_287_out;
    end
    endgenerate
    
    
    
    // LUT : 288
    wire [15:0] lut_288_table = 16'b1111001111110001;
    wire [3:0] lut_288_select = {
                             in_data[116],
                             in_data[277],
                             in_data[502],
                             in_data[273]};
    
    wire lut_288_out = lut_288_table[lut_288_select];
    
    generate
    if ( USE_REG ) begin : ff_288
        reg   lut_288_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_288_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_288_ff <= lut_288_out;
            end
        end
        
        assign out_data[288] = lut_288_ff;
    end
    else begin : no_ff_288
        assign out_data[288] = lut_288_out;
    end
    endgenerate
    
    
    
    // LUT : 289
    wire [15:0] lut_289_table = 16'b0100010101000100;
    wire [3:0] lut_289_select = {
                             in_data[211],
                             in_data[453],
                             in_data[68],
                             in_data[28]};
    
    wire lut_289_out = lut_289_table[lut_289_select];
    
    generate
    if ( USE_REG ) begin : ff_289
        reg   lut_289_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_289_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_289_ff <= lut_289_out;
            end
        end
        
        assign out_data[289] = lut_289_ff;
    end
    else begin : no_ff_289
        assign out_data[289] = lut_289_out;
    end
    endgenerate
    
    
    
    // LUT : 290
    wire [15:0] lut_290_table = 16'b0000110011001111;
    wire [3:0] lut_290_select = {
                             in_data[110],
                             in_data[234],
                             in_data[172],
                             in_data[213]};
    
    wire lut_290_out = lut_290_table[lut_290_select];
    
    generate
    if ( USE_REG ) begin : ff_290
        reg   lut_290_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_290_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_290_ff <= lut_290_out;
            end
        end
        
        assign out_data[290] = lut_290_ff;
    end
    else begin : no_ff_290
        assign out_data[290] = lut_290_out;
    end
    endgenerate
    
    
    
    // LUT : 291
    wire [15:0] lut_291_table = 16'b1010111110101110;
    wire [3:0] lut_291_select = {
                             in_data[170],
                             in_data[56],
                             in_data[494],
                             in_data[399]};
    
    wire lut_291_out = lut_291_table[lut_291_select];
    
    generate
    if ( USE_REG ) begin : ff_291
        reg   lut_291_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_291_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_291_ff <= lut_291_out;
            end
        end
        
        assign out_data[291] = lut_291_ff;
    end
    else begin : no_ff_291
        assign out_data[291] = lut_291_out;
    end
    endgenerate
    
    
    
    // LUT : 292
    wire [15:0] lut_292_table = 16'b0100010100000000;
    wire [3:0] lut_292_select = {
                             in_data[600],
                             in_data[311],
                             in_data[443],
                             in_data[47]};
    
    wire lut_292_out = lut_292_table[lut_292_select];
    
    generate
    if ( USE_REG ) begin : ff_292
        reg   lut_292_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_292_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_292_ff <= lut_292_out;
            end
        end
        
        assign out_data[292] = lut_292_ff;
    end
    else begin : no_ff_292
        assign out_data[292] = lut_292_out;
    end
    endgenerate
    
    
    
    // LUT : 293
    wire [15:0] lut_293_table = 16'b0000110011001100;
    wire [3:0] lut_293_select = {
                             in_data[214],
                             in_data[38],
                             in_data[636],
                             in_data[345]};
    
    wire lut_293_out = lut_293_table[lut_293_select];
    
    generate
    if ( USE_REG ) begin : ff_293
        reg   lut_293_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_293_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_293_ff <= lut_293_out;
            end
        end
        
        assign out_data[293] = lut_293_ff;
    end
    else begin : no_ff_293
        assign out_data[293] = lut_293_out;
    end
    endgenerate
    
    
    
    // LUT : 294
    wire [15:0] lut_294_table = 16'b1011000010110010;
    wire [3:0] lut_294_select = {
                             in_data[118],
                             in_data[274],
                             in_data[478],
                             in_data[250]};
    
    wire lut_294_out = lut_294_table[lut_294_select];
    
    generate
    if ( USE_REG ) begin : ff_294
        reg   lut_294_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_294_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_294_ff <= lut_294_out;
            end
        end
        
        assign out_data[294] = lut_294_ff;
    end
    else begin : no_ff_294
        assign out_data[294] = lut_294_out;
    end
    endgenerate
    
    
    
    // LUT : 295
    wire [15:0] lut_295_table = 16'b0000111100111111;
    wire [3:0] lut_295_select = {
                             in_data[469],
                             in_data[119],
                             in_data[483],
                             in_data[197]};
    
    wire lut_295_out = lut_295_table[lut_295_select];
    
    generate
    if ( USE_REG ) begin : ff_295
        reg   lut_295_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_295_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_295_ff <= lut_295_out;
            end
        end
        
        assign out_data[295] = lut_295_ff;
    end
    else begin : no_ff_295
        assign out_data[295] = lut_295_out;
    end
    endgenerate
    
    
    
    // LUT : 296
    wire [15:0] lut_296_table = 16'b0000010100000100;
    wire [3:0] lut_296_select = {
                             in_data[71],
                             in_data[135],
                             in_data[394],
                             in_data[182]};
    
    wire lut_296_out = lut_296_table[lut_296_select];
    
    generate
    if ( USE_REG ) begin : ff_296
        reg   lut_296_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_296_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_296_ff <= lut_296_out;
            end
        end
        
        assign out_data[296] = lut_296_ff;
    end
    else begin : no_ff_296
        assign out_data[296] = lut_296_out;
    end
    endgenerate
    
    
    
    // LUT : 297
    wire [15:0] lut_297_table = 16'b1010111100001010;
    wire [3:0] lut_297_select = {
                             in_data[330],
                             in_data[575],
                             in_data[507],
                             in_data[239]};
    
    wire lut_297_out = lut_297_table[lut_297_select];
    
    generate
    if ( USE_REG ) begin : ff_297
        reg   lut_297_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_297_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_297_ff <= lut_297_out;
            end
        end
        
        assign out_data[297] = lut_297_ff;
    end
    else begin : no_ff_297
        assign out_data[297] = lut_297_out;
    end
    endgenerate
    
    
    
    // LUT : 298
    wire [15:0] lut_298_table = 16'b1011101110111011;
    wire [3:0] lut_298_select = {
                             in_data[73],
                             in_data[329],
                             in_data[149],
                             in_data[422]};
    
    wire lut_298_out = lut_298_table[lut_298_select];
    
    generate
    if ( USE_REG ) begin : ff_298
        reg   lut_298_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_298_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_298_ff <= lut_298_out;
            end
        end
        
        assign out_data[298] = lut_298_ff;
    end
    else begin : no_ff_298
        assign out_data[298] = lut_298_out;
    end
    endgenerate
    
    
    
    // LUT : 299
    wire [15:0] lut_299_table = 16'b1011001100000011;
    wire [3:0] lut_299_select = {
                             in_data[573],
                             in_data[276],
                             in_data[433],
                             in_data[624]};
    
    wire lut_299_out = lut_299_table[lut_299_select];
    
    generate
    if ( USE_REG ) begin : ff_299
        reg   lut_299_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_299_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_299_ff <= lut_299_out;
            end
        end
        
        assign out_data[299] = lut_299_ff;
    end
    else begin : no_ff_299
        assign out_data[299] = lut_299_out;
    end
    endgenerate
    
    
    
    // LUT : 300
    wire [15:0] lut_300_table = 16'b1111111111110101;
    wire [3:0] lut_300_select = {
                             in_data[437],
                             in_data[594],
                             in_data[468],
                             in_data[263]};
    
    wire lut_300_out = lut_300_table[lut_300_select];
    
    generate
    if ( USE_REG ) begin : ff_300
        reg   lut_300_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_300_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_300_ff <= lut_300_out;
            end
        end
        
        assign out_data[300] = lut_300_ff;
    end
    else begin : no_ff_300
        assign out_data[300] = lut_300_out;
    end
    endgenerate
    
    
    
    // LUT : 301
    wire [15:0] lut_301_table = 16'b1010101011101000;
    wire [3:0] lut_301_select = {
                             in_data[360],
                             in_data[220],
                             in_data[142],
                             in_data[318]};
    
    wire lut_301_out = lut_301_table[lut_301_select];
    
    generate
    if ( USE_REG ) begin : ff_301
        reg   lut_301_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_301_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_301_ff <= lut_301_out;
            end
        end
        
        assign out_data[301] = lut_301_ff;
    end
    else begin : no_ff_301
        assign out_data[301] = lut_301_out;
    end
    endgenerate
    
    
    
    // LUT : 302
    wire [15:0] lut_302_table = 16'b0000000011111011;
    wire [3:0] lut_302_select = {
                             in_data[540],
                             in_data[432],
                             in_data[62],
                             in_data[34]};
    
    wire lut_302_out = lut_302_table[lut_302_select];
    
    generate
    if ( USE_REG ) begin : ff_302
        reg   lut_302_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_302_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_302_ff <= lut_302_out;
            end
        end
        
        assign out_data[302] = lut_302_ff;
    end
    else begin : no_ff_302
        assign out_data[302] = lut_302_out;
    end
    endgenerate
    
    
    
    // LUT : 303
    wire [15:0] lut_303_table = 16'b0000000000001111;
    wire [3:0] lut_303_select = {
                             in_data[417],
                             in_data[365],
                             in_data[459],
                             in_data[528]};
    
    wire lut_303_out = lut_303_table[lut_303_select];
    
    generate
    if ( USE_REG ) begin : ff_303
        reg   lut_303_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_303_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_303_ff <= lut_303_out;
            end
        end
        
        assign out_data[303] = lut_303_ff;
    end
    else begin : no_ff_303
        assign out_data[303] = lut_303_out;
    end
    endgenerate
    
    
    
    // LUT : 304
    wire [15:0] lut_304_table = 16'b1100000010101010;
    wire [3:0] lut_304_select = {
                             in_data[45],
                             in_data[532],
                             in_data[164],
                             in_data[50]};
    
    wire lut_304_out = lut_304_table[lut_304_select];
    
    generate
    if ( USE_REG ) begin : ff_304
        reg   lut_304_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_304_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_304_ff <= lut_304_out;
            end
        end
        
        assign out_data[304] = lut_304_ff;
    end
    else begin : no_ff_304
        assign out_data[304] = lut_304_out;
    end
    endgenerate
    
    
    
    // LUT : 305
    wire [15:0] lut_305_table = 16'b0001111100010111;
    wire [3:0] lut_305_select = {
                             in_data[307],
                             in_data[301],
                             in_data[114],
                             in_data[93]};
    
    wire lut_305_out = lut_305_table[lut_305_select];
    
    generate
    if ( USE_REG ) begin : ff_305
        reg   lut_305_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_305_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_305_ff <= lut_305_out;
            end
        end
        
        assign out_data[305] = lut_305_ff;
    end
    else begin : no_ff_305
        assign out_data[305] = lut_305_out;
    end
    endgenerate
    
    
    
    // LUT : 306
    wire [15:0] lut_306_table = 16'b0010111100000011;
    wire [3:0] lut_306_select = {
                             in_data[423],
                             in_data[166],
                             in_data[388],
                             in_data[27]};
    
    wire lut_306_out = lut_306_table[lut_306_select];
    
    generate
    if ( USE_REG ) begin : ff_306
        reg   lut_306_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_306_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_306_ff <= lut_306_out;
            end
        end
        
        assign out_data[306] = lut_306_ff;
    end
    else begin : no_ff_306
        assign out_data[306] = lut_306_out;
    end
    endgenerate
    
    
    
    // LUT : 307
    wire [15:0] lut_307_table = 16'b1011101100000000;
    wire [3:0] lut_307_select = {
                             in_data[84],
                             in_data[40],
                             in_data[403],
                             in_data[59]};
    
    wire lut_307_out = lut_307_table[lut_307_select];
    
    generate
    if ( USE_REG ) begin : ff_307
        reg   lut_307_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_307_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_307_ff <= lut_307_out;
            end
        end
        
        assign out_data[307] = lut_307_ff;
    end
    else begin : no_ff_307
        assign out_data[307] = lut_307_out;
    end
    endgenerate
    
    
    
    // LUT : 308
    wire [15:0] lut_308_table = 16'b0011001000110010;
    wire [3:0] lut_308_select = {
                             in_data[96],
                             in_data[463],
                             in_data[476],
                             in_data[209]};
    
    wire lut_308_out = lut_308_table[lut_308_select];
    
    generate
    if ( USE_REG ) begin : ff_308
        reg   lut_308_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_308_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_308_ff <= lut_308_out;
            end
        end
        
        assign out_data[308] = lut_308_ff;
    end
    else begin : no_ff_308
        assign out_data[308] = lut_308_out;
    end
    endgenerate
    
    
    
    // LUT : 309
    wire [15:0] lut_309_table = 16'b1111001111110011;
    wire [3:0] lut_309_select = {
                             in_data[635],
                             in_data[508],
                             in_data[639],
                             in_data[193]};
    
    wire lut_309_out = lut_309_table[lut_309_select];
    
    generate
    if ( USE_REG ) begin : ff_309
        reg   lut_309_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_309_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_309_ff <= lut_309_out;
            end
        end
        
        assign out_data[309] = lut_309_ff;
    end
    else begin : no_ff_309
        assign out_data[309] = lut_309_out;
    end
    endgenerate
    
    
    
    // LUT : 310
    wire [15:0] lut_310_table = 16'b1101010011010000;
    wire [3:0] lut_310_select = {
                             in_data[134],
                             in_data[103],
                             in_data[226],
                             in_data[613]};
    
    wire lut_310_out = lut_310_table[lut_310_select];
    
    generate
    if ( USE_REG ) begin : ff_310
        reg   lut_310_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_310_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_310_ff <= lut_310_out;
            end
        end
        
        assign out_data[310] = lut_310_ff;
    end
    else begin : no_ff_310
        assign out_data[310] = lut_310_out;
    end
    endgenerate
    
    
    
    // LUT : 311
    wire [15:0] lut_311_table = 16'b0000001101111111;
    wire [3:0] lut_311_select = {
                             in_data[121],
                             in_data[270],
                             in_data[570],
                             in_data[13]};
    
    wire lut_311_out = lut_311_table[lut_311_select];
    
    generate
    if ( USE_REG ) begin : ff_311
        reg   lut_311_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_311_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_311_ff <= lut_311_out;
            end
        end
        
        assign out_data[311] = lut_311_ff;
    end
    else begin : no_ff_311
        assign out_data[311] = lut_311_out;
    end
    endgenerate
    
    
    
    // LUT : 312
    wire [15:0] lut_312_table = 16'b1101111100000101;
    wire [3:0] lut_312_select = {
                             in_data[161],
                             in_data[3],
                             in_data[328],
                             in_data[288]};
    
    wire lut_312_out = lut_312_table[lut_312_select];
    
    generate
    if ( USE_REG ) begin : ff_312
        reg   lut_312_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_312_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_312_ff <= lut_312_out;
            end
        end
        
        assign out_data[312] = lut_312_ff;
    end
    else begin : no_ff_312
        assign out_data[312] = lut_312_out;
    end
    endgenerate
    
    
    
    // LUT : 313
    wire [15:0] lut_313_table = 16'b0101000000010000;
    wire [3:0] lut_313_select = {
                             in_data[499],
                             in_data[141],
                             in_data[362],
                             in_data[227]};
    
    wire lut_313_out = lut_313_table[lut_313_select];
    
    generate
    if ( USE_REG ) begin : ff_313
        reg   lut_313_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_313_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_313_ff <= lut_313_out;
            end
        end
        
        assign out_data[313] = lut_313_ff;
    end
    else begin : no_ff_313
        assign out_data[313] = lut_313_out;
    end
    endgenerate
    
    
    
    // LUT : 314
    wire [15:0] lut_314_table = 16'b1110111111001100;
    wire [3:0] lut_314_select = {
                             in_data[472],
                             in_data[560],
                             in_data[550],
                             in_data[136]};
    
    wire lut_314_out = lut_314_table[lut_314_select];
    
    generate
    if ( USE_REG ) begin : ff_314
        reg   lut_314_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_314_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_314_ff <= lut_314_out;
            end
        end
        
        assign out_data[314] = lut_314_ff;
    end
    else begin : no_ff_314
        assign out_data[314] = lut_314_out;
    end
    endgenerate
    
    
    
    // LUT : 315
    wire [15:0] lut_315_table = 16'b1111110011001100;
    wire [3:0] lut_315_select = {
                             in_data[597],
                             in_data[287],
                             in_data[279],
                             in_data[569]};
    
    wire lut_315_out = lut_315_table[lut_315_select];
    
    generate
    if ( USE_REG ) begin : ff_315
        reg   lut_315_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_315_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_315_ff <= lut_315_out;
            end
        end
        
        assign out_data[315] = lut_315_ff;
    end
    else begin : no_ff_315
        assign out_data[315] = lut_315_out;
    end
    endgenerate
    
    
    
    // LUT : 316
    wire [15:0] lut_316_table = 16'b0000001100001011;
    wire [3:0] lut_316_select = {
                             in_data[366],
                             in_data[336],
                             in_data[541],
                             in_data[420]};
    
    wire lut_316_out = lut_316_table[lut_316_select];
    
    generate
    if ( USE_REG ) begin : ff_316
        reg   lut_316_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_316_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_316_ff <= lut_316_out;
            end
        end
        
        assign out_data[316] = lut_316_ff;
    end
    else begin : no_ff_316
        assign out_data[316] = lut_316_out;
    end
    endgenerate
    
    
    
    // LUT : 317
    wire [15:0] lut_317_table = 16'b1111000011011000;
    wire [3:0] lut_317_select = {
                             in_data[405],
                             in_data[515],
                             in_data[292],
                             in_data[584]};
    
    wire lut_317_out = lut_317_table[lut_317_select];
    
    generate
    if ( USE_REG ) begin : ff_317
        reg   lut_317_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_317_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_317_ff <= lut_317_out;
            end
        end
        
        assign out_data[317] = lut_317_ff;
    end
    else begin : no_ff_317
        assign out_data[317] = lut_317_out;
    end
    endgenerate
    
    
    
    // LUT : 318
    wire [15:0] lut_318_table = 16'b0011001111110011;
    wire [3:0] lut_318_select = {
                             in_data[87],
                             in_data[58],
                             in_data[421],
                             in_data[340]};
    
    wire lut_318_out = lut_318_table[lut_318_select];
    
    generate
    if ( USE_REG ) begin : ff_318
        reg   lut_318_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_318_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_318_ff <= lut_318_out;
            end
        end
        
        assign out_data[318] = lut_318_ff;
    end
    else begin : no_ff_318
        assign out_data[318] = lut_318_out;
    end
    endgenerate
    
    
    
    // LUT : 319
    wire [15:0] lut_319_table = 16'b0111000111110001;
    wire [3:0] lut_319_select = {
                             in_data[375],
                             in_data[207],
                             in_data[251],
                             in_data[390]};
    
    wire lut_319_out = lut_319_table[lut_319_select];
    
    generate
    if ( USE_REG ) begin : ff_319
        reg   lut_319_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_319_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_319_ff <= lut_319_out;
            end
        end
        
        assign out_data[319] = lut_319_ff;
    end
    else begin : no_ff_319
        assign out_data[319] = lut_319_out;
    end
    endgenerate
    
    
    
    // LUT : 320
    wire [15:0] lut_320_table = 16'b0000000101010111;
    wire [3:0] lut_320_select = {
                             in_data[615],
                             in_data[366],
                             in_data[52],
                             in_data[235]};
    
    wire lut_320_out = lut_320_table[lut_320_select];
    
    generate
    if ( USE_REG ) begin : ff_320
        reg   lut_320_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_320_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_320_ff <= lut_320_out;
            end
        end
        
        assign out_data[320] = lut_320_ff;
    end
    else begin : no_ff_320
        assign out_data[320] = lut_320_out;
    end
    endgenerate
    
    
    
    // LUT : 321
    wire [15:0] lut_321_table = 16'b0001000111110111;
    wire [3:0] lut_321_select = {
                             in_data[477],
                             in_data[561],
                             in_data[273],
                             in_data[291]};
    
    wire lut_321_out = lut_321_table[lut_321_select];
    
    generate
    if ( USE_REG ) begin : ff_321
        reg   lut_321_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_321_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_321_ff <= lut_321_out;
            end
        end
        
        assign out_data[321] = lut_321_ff;
    end
    else begin : no_ff_321
        assign out_data[321] = lut_321_out;
    end
    endgenerate
    
    
    
    // LUT : 322
    wire [15:0] lut_322_table = 16'b0000000100110011;
    wire [3:0] lut_322_select = {
                             in_data[468],
                             in_data[338],
                             in_data[219],
                             in_data[451]};
    
    wire lut_322_out = lut_322_table[lut_322_select];
    
    generate
    if ( USE_REG ) begin : ff_322
        reg   lut_322_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_322_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_322_ff <= lut_322_out;
            end
        end
        
        assign out_data[322] = lut_322_ff;
    end
    else begin : no_ff_322
        assign out_data[322] = lut_322_out;
    end
    endgenerate
    
    
    
    // LUT : 323
    wire [15:0] lut_323_table = 16'b1111111100000111;
    wire [3:0] lut_323_select = {
                             in_data[70],
                             in_data[398],
                             in_data[414],
                             in_data[147]};
    
    wire lut_323_out = lut_323_table[lut_323_select];
    
    generate
    if ( USE_REG ) begin : ff_323
        reg   lut_323_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_323_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_323_ff <= lut_323_out;
            end
        end
        
        assign out_data[323] = lut_323_ff;
    end
    else begin : no_ff_323
        assign out_data[323] = lut_323_out;
    end
    endgenerate
    
    
    
    // LUT : 324
    wire [15:0] lut_324_table = 16'b1111111100001111;
    wire [3:0] lut_324_select = {
                             in_data[552],
                             in_data[153],
                             in_data[631],
                             in_data[108]};
    
    wire lut_324_out = lut_324_table[lut_324_select];
    
    generate
    if ( USE_REG ) begin : ff_324
        reg   lut_324_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_324_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_324_ff <= lut_324_out;
            end
        end
        
        assign out_data[324] = lut_324_ff;
    end
    else begin : no_ff_324
        assign out_data[324] = lut_324_out;
    end
    endgenerate
    
    
    
    // LUT : 325
    wire [15:0] lut_325_table = 16'b1010000011110001;
    wire [3:0] lut_325_select = {
                             in_data[349],
                             in_data[433],
                             in_data[154],
                             in_data[324]};
    
    wire lut_325_out = lut_325_table[lut_325_select];
    
    generate
    if ( USE_REG ) begin : ff_325
        reg   lut_325_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_325_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_325_ff <= lut_325_out;
            end
        end
        
        assign out_data[325] = lut_325_ff;
    end
    else begin : no_ff_325
        assign out_data[325] = lut_325_out;
    end
    endgenerate
    
    
    
    // LUT : 326
    wire [15:0] lut_326_table = 16'b0101010011110101;
    wire [3:0] lut_326_select = {
                             in_data[55],
                             in_data[21],
                             in_data[590],
                             in_data[353]};
    
    wire lut_326_out = lut_326_table[lut_326_select];
    
    generate
    if ( USE_REG ) begin : ff_326
        reg   lut_326_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_326_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_326_ff <= lut_326_out;
            end
        end
        
        assign out_data[326] = lut_326_ff;
    end
    else begin : no_ff_326
        assign out_data[326] = lut_326_out;
    end
    endgenerate
    
    
    
    // LUT : 327
    wire [15:0] lut_327_table = 16'b0000100010101110;
    wire [3:0] lut_327_select = {
                             in_data[286],
                             in_data[604],
                             in_data[464],
                             in_data[405]};
    
    wire lut_327_out = lut_327_table[lut_327_select];
    
    generate
    if ( USE_REG ) begin : ff_327
        reg   lut_327_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_327_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_327_ff <= lut_327_out;
            end
        end
        
        assign out_data[327] = lut_327_ff;
    end
    else begin : no_ff_327
        assign out_data[327] = lut_327_out;
    end
    endgenerate
    
    
    
    // LUT : 328
    wire [15:0] lut_328_table = 16'b0000000011101100;
    wire [3:0] lut_328_select = {
                             in_data[429],
                             in_data[35],
                             in_data[133],
                             in_data[438]};
    
    wire lut_328_out = lut_328_table[lut_328_select];
    
    generate
    if ( USE_REG ) begin : ff_328
        reg   lut_328_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_328_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_328_ff <= lut_328_out;
            end
        end
        
        assign out_data[328] = lut_328_ff;
    end
    else begin : no_ff_328
        assign out_data[328] = lut_328_out;
    end
    endgenerate
    
    
    
    // LUT : 329
    wire [15:0] lut_329_table = 16'b0000000000001111;
    wire [3:0] lut_329_select = {
                             in_data[471],
                             in_data[166],
                             in_data[305],
                             in_data[387]};
    
    wire lut_329_out = lut_329_table[lut_329_select];
    
    generate
    if ( USE_REG ) begin : ff_329
        reg   lut_329_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_329_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_329_ff <= lut_329_out;
            end
        end
        
        assign out_data[329] = lut_329_ff;
    end
    else begin : no_ff_329
        assign out_data[329] = lut_329_out;
    end
    endgenerate
    
    
    
    // LUT : 330
    wire [15:0] lut_330_table = 16'b1000100010001000;
    wire [3:0] lut_330_select = {
                             in_data[453],
                             in_data[634],
                             in_data[90],
                             in_data[8]};
    
    wire lut_330_out = lut_330_table[lut_330_select];
    
    generate
    if ( USE_REG ) begin : ff_330
        reg   lut_330_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_330_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_330_ff <= lut_330_out;
            end
        end
        
        assign out_data[330] = lut_330_ff;
    end
    else begin : no_ff_330
        assign out_data[330] = lut_330_out;
    end
    endgenerate
    
    
    
    // LUT : 331
    wire [15:0] lut_331_table = 16'b0101110001011101;
    wire [3:0] lut_331_select = {
                             in_data[180],
                             in_data[268],
                             in_data[174],
                             in_data[51]};
    
    wire lut_331_out = lut_331_table[lut_331_select];
    
    generate
    if ( USE_REG ) begin : ff_331
        reg   lut_331_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_331_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_331_ff <= lut_331_out;
            end
        end
        
        assign out_data[331] = lut_331_ff;
    end
    else begin : no_ff_331
        assign out_data[331] = lut_331_out;
    end
    endgenerate
    
    
    
    // LUT : 332
    wire [15:0] lut_332_table = 16'b1100110011001100;
    wire [3:0] lut_332_select = {
                             in_data[53],
                             in_data[261],
                             in_data[298],
                             in_data[56]};
    
    wire lut_332_out = lut_332_table[lut_332_select];
    
    generate
    if ( USE_REG ) begin : ff_332
        reg   lut_332_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_332_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_332_ff <= lut_332_out;
            end
        end
        
        assign out_data[332] = lut_332_ff;
    end
    else begin : no_ff_332
        assign out_data[332] = lut_332_out;
    end
    endgenerate
    
    
    
    // LUT : 333
    wire [15:0] lut_333_table = 16'b1110110011101100;
    wire [3:0] lut_333_select = {
                             in_data[524],
                             in_data[170],
                             in_data[132],
                             in_data[284]};
    
    wire lut_333_out = lut_333_table[lut_333_select];
    
    generate
    if ( USE_REG ) begin : ff_333
        reg   lut_333_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_333_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_333_ff <= lut_333_out;
            end
        end
        
        assign out_data[333] = lut_333_ff;
    end
    else begin : no_ff_333
        assign out_data[333] = lut_333_out;
    end
    endgenerate
    
    
    
    // LUT : 334
    wire [15:0] lut_334_table = 16'b0100111011001111;
    wire [3:0] lut_334_select = {
                             in_data[421],
                             in_data[584],
                             in_data[345],
                             in_data[500]};
    
    wire lut_334_out = lut_334_table[lut_334_select];
    
    generate
    if ( USE_REG ) begin : ff_334
        reg   lut_334_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_334_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_334_ff <= lut_334_out;
            end
        end
        
        assign out_data[334] = lut_334_ff;
    end
    else begin : no_ff_334
        assign out_data[334] = lut_334_out;
    end
    endgenerate
    
    
    
    // LUT : 335
    wire [15:0] lut_335_table = 16'b0111000111110000;
    wire [3:0] lut_335_select = {
                             in_data[136],
                             in_data[206],
                             in_data[44],
                             in_data[274]};
    
    wire lut_335_out = lut_335_table[lut_335_select];
    
    generate
    if ( USE_REG ) begin : ff_335
        reg   lut_335_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_335_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_335_ff <= lut_335_out;
            end
        end
        
        assign out_data[335] = lut_335_ff;
    end
    else begin : no_ff_335
        assign out_data[335] = lut_335_out;
    end
    endgenerate
    
    
    
    // LUT : 336
    wire [15:0] lut_336_table = 16'b1111101011111010;
    wire [3:0] lut_336_select = {
                             in_data[550],
                             in_data[517],
                             in_data[49],
                             in_data[583]};
    
    wire lut_336_out = lut_336_table[lut_336_select];
    
    generate
    if ( USE_REG ) begin : ff_336
        reg   lut_336_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_336_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_336_ff <= lut_336_out;
            end
        end
        
        assign out_data[336] = lut_336_ff;
    end
    else begin : no_ff_336
        assign out_data[336] = lut_336_out;
    end
    endgenerate
    
    
    
    // LUT : 337
    wire [15:0] lut_337_table = 16'b0100010100000101;
    wire [3:0] lut_337_select = {
                             in_data[97],
                             in_data[603],
                             in_data[490],
                             in_data[367]};
    
    wire lut_337_out = lut_337_table[lut_337_select];
    
    generate
    if ( USE_REG ) begin : ff_337
        reg   lut_337_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_337_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_337_ff <= lut_337_out;
            end
        end
        
        assign out_data[337] = lut_337_ff;
    end
    else begin : no_ff_337
        assign out_data[337] = lut_337_out;
    end
    endgenerate
    
    
    
    // LUT : 338
    wire [15:0] lut_338_table = 16'b0101000101010001;
    wire [3:0] lut_338_select = {
                             in_data[62],
                             in_data[492],
                             in_data[466],
                             in_data[611]};
    
    wire lut_338_out = lut_338_table[lut_338_select];
    
    generate
    if ( USE_REG ) begin : ff_338
        reg   lut_338_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_338_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_338_ff <= lut_338_out;
            end
        end
        
        assign out_data[338] = lut_338_ff;
    end
    else begin : no_ff_338
        assign out_data[338] = lut_338_out;
    end
    endgenerate
    
    
    
    // LUT : 339
    wire [15:0] lut_339_table = 16'b1111111011111100;
    wire [3:0] lut_339_select = {
                             in_data[616],
                             in_data[225],
                             in_data[446],
                             in_data[276]};
    
    wire lut_339_out = lut_339_table[lut_339_select];
    
    generate
    if ( USE_REG ) begin : ff_339
        reg   lut_339_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_339_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_339_ff <= lut_339_out;
            end
        end
        
        assign out_data[339] = lut_339_ff;
    end
    else begin : no_ff_339
        assign out_data[339] = lut_339_out;
    end
    endgenerate
    
    
    
    // LUT : 340
    wire [15:0] lut_340_table = 16'b0101010101000101;
    wire [3:0] lut_340_select = {
                             in_data[80],
                             in_data[407],
                             in_data[502],
                             in_data[327]};
    
    wire lut_340_out = lut_340_table[lut_340_select];
    
    generate
    if ( USE_REG ) begin : ff_340
        reg   lut_340_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_340_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_340_ff <= lut_340_out;
            end
        end
        
        assign out_data[340] = lut_340_ff;
    end
    else begin : no_ff_340
        assign out_data[340] = lut_340_out;
    end
    endgenerate
    
    
    
    // LUT : 341
    wire [15:0] lut_341_table = 16'b1111011100110011;
    wire [3:0] lut_341_select = {
                             in_data[242],
                             in_data[119],
                             in_data[110],
                             in_data[222]};
    
    wire lut_341_out = lut_341_table[lut_341_select];
    
    generate
    if ( USE_REG ) begin : ff_341
        reg   lut_341_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_341_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_341_ff <= lut_341_out;
            end
        end
        
        assign out_data[341] = lut_341_ff;
    end
    else begin : no_ff_341
        assign out_data[341] = lut_341_out;
    end
    endgenerate
    
    
    
    // LUT : 342
    wire [15:0] lut_342_table = 16'b0000000011101111;
    wire [3:0] lut_342_select = {
                             in_data[486],
                             in_data[200],
                             in_data[636],
                             in_data[272]};
    
    wire lut_342_out = lut_342_table[lut_342_select];
    
    generate
    if ( USE_REG ) begin : ff_342
        reg   lut_342_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_342_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_342_ff <= lut_342_out;
            end
        end
        
        assign out_data[342] = lut_342_ff;
    end
    else begin : no_ff_342
        assign out_data[342] = lut_342_out;
    end
    endgenerate
    
    
    
    // LUT : 343
    wire [15:0] lut_343_table = 16'b0000111100000010;
    wire [3:0] lut_343_select = {
                             in_data[211],
                             in_data[168],
                             in_data[411],
                             in_data[114]};
    
    wire lut_343_out = lut_343_table[lut_343_select];
    
    generate
    if ( USE_REG ) begin : ff_343
        reg   lut_343_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_343_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_343_ff <= lut_343_out;
            end
        end
        
        assign out_data[343] = lut_343_ff;
    end
    else begin : no_ff_343
        assign out_data[343] = lut_343_out;
    end
    endgenerate
    
    
    
    // LUT : 344
    wire [15:0] lut_344_table = 16'b1111100011110000;
    wire [3:0] lut_344_select = {
                             in_data[428],
                             in_data[511],
                             in_data[248],
                             in_data[107]};
    
    wire lut_344_out = lut_344_table[lut_344_select];
    
    generate
    if ( USE_REG ) begin : ff_344
        reg   lut_344_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_344_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_344_ff <= lut_344_out;
            end
        end
        
        assign out_data[344] = lut_344_ff;
    end
    else begin : no_ff_344
        assign out_data[344] = lut_344_out;
    end
    endgenerate
    
    
    
    // LUT : 345
    wire [15:0] lut_345_table = 16'b1111010011000100;
    wire [3:0] lut_345_select = {
                             in_data[176],
                             in_data[165],
                             in_data[295],
                             in_data[385]};
    
    wire lut_345_out = lut_345_table[lut_345_select];
    
    generate
    if ( USE_REG ) begin : ff_345
        reg   lut_345_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_345_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_345_ff <= lut_345_out;
            end
        end
        
        assign out_data[345] = lut_345_ff;
    end
    else begin : no_ff_345
        assign out_data[345] = lut_345_out;
    end
    endgenerate
    
    
    
    // LUT : 346
    wire [15:0] lut_346_table = 16'b1111110111011100;
    wire [3:0] lut_346_select = {
                             in_data[104],
                             in_data[263],
                             in_data[410],
                             in_data[0]};
    
    wire lut_346_out = lut_346_table[lut_346_select];
    
    generate
    if ( USE_REG ) begin : ff_346
        reg   lut_346_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_346_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_346_ff <= lut_346_out;
            end
        end
        
        assign out_data[346] = lut_346_ff;
    end
    else begin : no_ff_346
        assign out_data[346] = lut_346_out;
    end
    endgenerate
    
    
    
    // LUT : 347
    wire [15:0] lut_347_table = 16'b1111010011110000;
    wire [3:0] lut_347_select = {
                             in_data[621],
                             in_data[565],
                             in_data[279],
                             in_data[356]};
    
    wire lut_347_out = lut_347_table[lut_347_select];
    
    generate
    if ( USE_REG ) begin : ff_347
        reg   lut_347_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_347_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_347_ff <= lut_347_out;
            end
        end
        
        assign out_data[347] = lut_347_ff;
    end
    else begin : no_ff_347
        assign out_data[347] = lut_347_out;
    end
    endgenerate
    
    
    
    // LUT : 348
    wire [15:0] lut_348_table = 16'b0100111100000000;
    wire [3:0] lut_348_select = {
                             in_data[193],
                             in_data[521],
                             in_data[149],
                             in_data[11]};
    
    wire lut_348_out = lut_348_table[lut_348_select];
    
    generate
    if ( USE_REG ) begin : ff_348
        reg   lut_348_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_348_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_348_ff <= lut_348_out;
            end
        end
        
        assign out_data[348] = lut_348_ff;
    end
    else begin : no_ff_348
        assign out_data[348] = lut_348_out;
    end
    endgenerate
    
    
    
    // LUT : 349
    wire [15:0] lut_349_table = 16'b0010000000101010;
    wire [3:0] lut_349_select = {
                             in_data[232],
                             in_data[607],
                             in_data[637],
                             in_data[573]};
    
    wire lut_349_out = lut_349_table[lut_349_select];
    
    generate
    if ( USE_REG ) begin : ff_349
        reg   lut_349_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_349_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_349_ff <= lut_349_out;
            end
        end
        
        assign out_data[349] = lut_349_ff;
    end
    else begin : no_ff_349
        assign out_data[349] = lut_349_out;
    end
    endgenerate
    
    
    
    // LUT : 350
    wire [15:0] lut_350_table = 16'b0100000001010100;
    wire [3:0] lut_350_select = {
                             in_data[626],
                             in_data[37],
                             in_data[638],
                             in_data[60]};
    
    wire lut_350_out = lut_350_table[lut_350_select];
    
    generate
    if ( USE_REG ) begin : ff_350
        reg   lut_350_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_350_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_350_ff <= lut_350_out;
            end
        end
        
        assign out_data[350] = lut_350_ff;
    end
    else begin : no_ff_350
        assign out_data[350] = lut_350_out;
    end
    endgenerate
    
    
    
    // LUT : 351
    wire [15:0] lut_351_table = 16'b1111011101010001;
    wire [3:0] lut_351_select = {
                             in_data[150],
                             in_data[197],
                             in_data[533],
                             in_data[333]};
    
    wire lut_351_out = lut_351_table[lut_351_select];
    
    generate
    if ( USE_REG ) begin : ff_351
        reg   lut_351_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_351_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_351_ff <= lut_351_out;
            end
        end
        
        assign out_data[351] = lut_351_ff;
    end
    else begin : no_ff_351
        assign out_data[351] = lut_351_out;
    end
    endgenerate
    
    
    
    // LUT : 352
    wire [15:0] lut_352_table = 16'b0111001100010001;
    wire [3:0] lut_352_select = {
                             in_data[258],
                             in_data[39],
                             in_data[138],
                             in_data[98]};
    
    wire lut_352_out = lut_352_table[lut_352_select];
    
    generate
    if ( USE_REG ) begin : ff_352
        reg   lut_352_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_352_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_352_ff <= lut_352_out;
            end
        end
        
        assign out_data[352] = lut_352_ff;
    end
    else begin : no_ff_352
        assign out_data[352] = lut_352_out;
    end
    endgenerate
    
    
    
    // LUT : 353
    wire [15:0] lut_353_table = 16'b0111011101110111;
    wire [3:0] lut_353_select = {
                             in_data[31],
                             in_data[280],
                             in_data[470],
                             in_data[74]};
    
    wire lut_353_out = lut_353_table[lut_353_select];
    
    generate
    if ( USE_REG ) begin : ff_353
        reg   lut_353_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_353_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_353_ff <= lut_353_out;
            end
        end
        
        assign out_data[353] = lut_353_ff;
    end
    else begin : no_ff_353
        assign out_data[353] = lut_353_out;
    end
    endgenerate
    
    
    
    // LUT : 354
    wire [15:0] lut_354_table = 16'b0111101100010000;
    wire [3:0] lut_354_select = {
                             in_data[59],
                             in_data[518],
                             in_data[192],
                             in_data[159]};
    
    wire lut_354_out = lut_354_table[lut_354_select];
    
    generate
    if ( USE_REG ) begin : ff_354
        reg   lut_354_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_354_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_354_ff <= lut_354_out;
            end
        end
        
        assign out_data[354] = lut_354_ff;
    end
    else begin : no_ff_354
        assign out_data[354] = lut_354_out;
    end
    endgenerate
    
    
    
    // LUT : 355
    wire [15:0] lut_355_table = 16'b0000111100100111;
    wire [3:0] lut_355_select = {
                             in_data[337],
                             in_data[188],
                             in_data[121],
                             in_data[409]};
    
    wire lut_355_out = lut_355_table[lut_355_select];
    
    generate
    if ( USE_REG ) begin : ff_355
        reg   lut_355_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_355_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_355_ff <= lut_355_out;
            end
        end
        
        assign out_data[355] = lut_355_ff;
    end
    else begin : no_ff_355
        assign out_data[355] = lut_355_out;
    end
    endgenerate
    
    
    
    // LUT : 356
    wire [15:0] lut_356_table = 16'b1100000011010100;
    wire [3:0] lut_356_select = {
                             in_data[122],
                             in_data[5],
                             in_data[13],
                             in_data[294]};
    
    wire lut_356_out = lut_356_table[lut_356_select];
    
    generate
    if ( USE_REG ) begin : ff_356
        reg   lut_356_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_356_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_356_ff <= lut_356_out;
            end
        end
        
        assign out_data[356] = lut_356_ff;
    end
    else begin : no_ff_356
        assign out_data[356] = lut_356_out;
    end
    endgenerate
    
    
    
    // LUT : 357
    wire [15:0] lut_357_table = 16'b0101010100000000;
    wire [3:0] lut_357_select = {
                             in_data[113],
                             in_data[506],
                             in_data[134],
                             in_data[450]};
    
    wire lut_357_out = lut_357_table[lut_357_select];
    
    generate
    if ( USE_REG ) begin : ff_357
        reg   lut_357_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_357_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_357_ff <= lut_357_out;
            end
        end
        
        assign out_data[357] = lut_357_ff;
    end
    else begin : no_ff_357
        assign out_data[357] = lut_357_out;
    end
    endgenerate
    
    
    
    // LUT : 358
    wire [15:0] lut_358_table = 16'b1111111111011100;
    wire [3:0] lut_358_select = {
                             in_data[162],
                             in_data[539],
                             in_data[260],
                             in_data[443]};
    
    wire lut_358_out = lut_358_table[lut_358_select];
    
    generate
    if ( USE_REG ) begin : ff_358
        reg   lut_358_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_358_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_358_ff <= lut_358_out;
            end
        end
        
        assign out_data[358] = lut_358_ff;
    end
    else begin : no_ff_358
        assign out_data[358] = lut_358_out;
    end
    endgenerate
    
    
    
    // LUT : 359
    wire [15:0] lut_359_table = 16'b0000000010111001;
    wire [3:0] lut_359_select = {
                             in_data[633],
                             in_data[448],
                             in_data[553],
                             in_data[283]};
    
    wire lut_359_out = lut_359_table[lut_359_select];
    
    generate
    if ( USE_REG ) begin : ff_359
        reg   lut_359_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_359_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_359_ff <= lut_359_out;
            end
        end
        
        assign out_data[359] = lut_359_ff;
    end
    else begin : no_ff_359
        assign out_data[359] = lut_359_out;
    end
    endgenerate
    
    
    
    // LUT : 360
    wire [15:0] lut_360_table = 16'b1010101100101010;
    wire [3:0] lut_360_select = {
                             in_data[36],
                             in_data[529],
                             in_data[83],
                             in_data[308]};
    
    wire lut_360_out = lut_360_table[lut_360_select];
    
    generate
    if ( USE_REG ) begin : ff_360
        reg   lut_360_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_360_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_360_ff <= lut_360_out;
            end
        end
        
        assign out_data[360] = lut_360_ff;
    end
    else begin : no_ff_360
        assign out_data[360] = lut_360_out;
    end
    endgenerate
    
    
    
    // LUT : 361
    wire [15:0] lut_361_table = 16'b1011111110101110;
    wire [3:0] lut_361_select = {
                             in_data[190],
                             in_data[544],
                             in_data[579],
                             in_data[434]};
    
    wire lut_361_out = lut_361_table[lut_361_select];
    
    generate
    if ( USE_REG ) begin : ff_361
        reg   lut_361_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_361_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_361_ff <= lut_361_out;
            end
        end
        
        assign out_data[361] = lut_361_ff;
    end
    else begin : no_ff_361
        assign out_data[361] = lut_361_out;
    end
    endgenerate
    
    
    
    // LUT : 362
    wire [15:0] lut_362_table = 16'b0000010101001101;
    wire [3:0] lut_362_select = {
                             in_data[16],
                             in_data[538],
                             in_data[447],
                             in_data[473]};
    
    wire lut_362_out = lut_362_table[lut_362_select];
    
    generate
    if ( USE_REG ) begin : ff_362
        reg   lut_362_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_362_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_362_ff <= lut_362_out;
            end
        end
        
        assign out_data[362] = lut_362_ff;
    end
    else begin : no_ff_362
        assign out_data[362] = lut_362_out;
    end
    endgenerate
    
    
    
    // LUT : 363
    wire [15:0] lut_363_table = 16'b1010101000000000;
    wire [3:0] lut_363_select = {
                             in_data[632],
                             in_data[559],
                             in_data[230],
                             in_data[396]};
    
    wire lut_363_out = lut_363_table[lut_363_select];
    
    generate
    if ( USE_REG ) begin : ff_363
        reg   lut_363_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_363_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_363_ff <= lut_363_out;
            end
        end
        
        assign out_data[363] = lut_363_ff;
    end
    else begin : no_ff_363
        assign out_data[363] = lut_363_out;
    end
    endgenerate
    
    
    
    // LUT : 364
    wire [15:0] lut_364_table = 16'b1111101011110010;
    wire [3:0] lut_364_select = {
                             in_data[600],
                             in_data[493],
                             in_data[487],
                             in_data[424]};
    
    wire lut_364_out = lut_364_table[lut_364_select];
    
    generate
    if ( USE_REG ) begin : ff_364
        reg   lut_364_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_364_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_364_ff <= lut_364_out;
            end
        end
        
        assign out_data[364] = lut_364_ff;
    end
    else begin : no_ff_364
        assign out_data[364] = lut_364_out;
    end
    endgenerate
    
    
    
    // LUT : 365
    wire [15:0] lut_365_table = 16'b1000000011111100;
    wire [3:0] lut_365_select = {
                             in_data[478],
                             in_data[588],
                             in_data[381],
                             in_data[129]};
    
    wire lut_365_out = lut_365_table[lut_365_select];
    
    generate
    if ( USE_REG ) begin : ff_365
        reg   lut_365_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_365_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_365_ff <= lut_365_out;
            end
        end
        
        assign out_data[365] = lut_365_ff;
    end
    else begin : no_ff_365
        assign out_data[365] = lut_365_out;
    end
    endgenerate
    
    
    
    // LUT : 366
    wire [15:0] lut_366_table = 16'b1111010101110101;
    wire [3:0] lut_366_select = {
                             in_data[370],
                             in_data[25],
                             in_data[629],
                             in_data[292]};
    
    wire lut_366_out = lut_366_table[lut_366_select];
    
    generate
    if ( USE_REG ) begin : ff_366
        reg   lut_366_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_366_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_366_ff <= lut_366_out;
            end
        end
        
        assign out_data[366] = lut_366_ff;
    end
    else begin : no_ff_366
        assign out_data[366] = lut_366_out;
    end
    endgenerate
    
    
    
    // LUT : 367
    wire [15:0] lut_367_table = 16'b1111101010100000;
    wire [3:0] lut_367_select = {
                             in_data[93],
                             in_data[256],
                             in_data[560],
                             in_data[392]};
    
    wire lut_367_out = lut_367_table[lut_367_select];
    
    generate
    if ( USE_REG ) begin : ff_367
        reg   lut_367_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_367_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_367_ff <= lut_367_out;
            end
        end
        
        assign out_data[367] = lut_367_ff;
    end
    else begin : no_ff_367
        assign out_data[367] = lut_367_out;
    end
    endgenerate
    
    
    
    // LUT : 368
    wire [15:0] lut_368_table = 16'b0101010101111111;
    wire [3:0] lut_368_select = {
                             in_data[509],
                             in_data[397],
                             in_data[460],
                             in_data[40]};
    
    wire lut_368_out = lut_368_table[lut_368_select];
    
    generate
    if ( USE_REG ) begin : ff_368
        reg   lut_368_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_368_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_368_ff <= lut_368_out;
            end
        end
        
        assign out_data[368] = lut_368_ff;
    end
    else begin : no_ff_368
        assign out_data[368] = lut_368_out;
    end
    endgenerate
    
    
    
    // LUT : 369
    wire [15:0] lut_369_table = 16'b0000010101111111;
    wire [3:0] lut_369_select = {
                             in_data[505],
                             in_data[599],
                             in_data[557],
                             in_data[362]};
    
    wire lut_369_out = lut_369_table[lut_369_select];
    
    generate
    if ( USE_REG ) begin : ff_369
        reg   lut_369_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_369_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_369_ff <= lut_369_out;
            end
        end
        
        assign out_data[369] = lut_369_ff;
    end
    else begin : no_ff_369
        assign out_data[369] = lut_369_out;
    end
    endgenerate
    
    
    
    // LUT : 370
    wire [15:0] lut_370_table = 16'b1010100011101010;
    wire [3:0] lut_370_select = {
                             in_data[281],
                             in_data[365],
                             in_data[204],
                             in_data[311]};
    
    wire lut_370_out = lut_370_table[lut_370_select];
    
    generate
    if ( USE_REG ) begin : ff_370
        reg   lut_370_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_370_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_370_ff <= lut_370_out;
            end
        end
        
        assign out_data[370] = lut_370_ff;
    end
    else begin : no_ff_370
        assign out_data[370] = lut_370_out;
    end
    endgenerate
    
    
    
    // LUT : 371
    wire [15:0] lut_371_table = 16'b0011111100000000;
    wire [3:0] lut_371_select = {
                             in_data[580],
                             in_data[540],
                             in_data[419],
                             in_data[507]};
    
    wire lut_371_out = lut_371_table[lut_371_select];
    
    generate
    if ( USE_REG ) begin : ff_371
        reg   lut_371_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_371_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_371_ff <= lut_371_out;
            end
        end
        
        assign out_data[371] = lut_371_ff;
    end
    else begin : no_ff_371
        assign out_data[371] = lut_371_out;
    end
    endgenerate
    
    
    
    // LUT : 372
    wire [15:0] lut_372_table = 16'b0000000011111111;
    wire [3:0] lut_372_select = {
                             in_data[253],
                             in_data[306],
                             in_data[569],
                             in_data[556]};
    
    wire lut_372_out = lut_372_table[lut_372_select];
    
    generate
    if ( USE_REG ) begin : ff_372
        reg   lut_372_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_372_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_372_ff <= lut_372_out;
            end
        end
        
        assign out_data[372] = lut_372_ff;
    end
    else begin : no_ff_372
        assign out_data[372] = lut_372_out;
    end
    endgenerate
    
    
    
    // LUT : 373
    wire [15:0] lut_373_table = 16'b1101010001000000;
    wire [3:0] lut_373_select = {
                             in_data[564],
                             in_data[151],
                             in_data[304],
                             in_data[426]};
    
    wire lut_373_out = lut_373_table[lut_373_select];
    
    generate
    if ( USE_REG ) begin : ff_373
        reg   lut_373_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_373_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_373_ff <= lut_373_out;
            end
        end
        
        assign out_data[373] = lut_373_ff;
    end
    else begin : no_ff_373
        assign out_data[373] = lut_373_out;
    end
    endgenerate
    
    
    
    // LUT : 374
    wire [15:0] lut_374_table = 16'b1101110111000100;
    wire [3:0] lut_374_select = {
                             in_data[47],
                             in_data[329],
                             in_data[30],
                             in_data[578]};
    
    wire lut_374_out = lut_374_table[lut_374_select];
    
    generate
    if ( USE_REG ) begin : ff_374
        reg   lut_374_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_374_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_374_ff <= lut_374_out;
            end
        end
        
        assign out_data[374] = lut_374_ff;
    end
    else begin : no_ff_374
        assign out_data[374] = lut_374_out;
    end
    endgenerate
    
    
    
    // LUT : 375
    wire [15:0] lut_375_table = 16'b0011001100110011;
    wire [3:0] lut_375_select = {
                             in_data[610],
                             in_data[591],
                             in_data[6],
                             in_data[315]};
    
    wire lut_375_out = lut_375_table[lut_375_select];
    
    generate
    if ( USE_REG ) begin : ff_375
        reg   lut_375_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_375_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_375_ff <= lut_375_out;
            end
        end
        
        assign out_data[375] = lut_375_ff;
    end
    else begin : no_ff_375
        assign out_data[375] = lut_375_out;
    end
    endgenerate
    
    
    
    // LUT : 376
    wire [15:0] lut_376_table = 16'b0000011100000000;
    wire [3:0] lut_376_select = {
                             in_data[501],
                             in_data[290],
                             in_data[627],
                             in_data[449]};
    
    wire lut_376_out = lut_376_table[lut_376_select];
    
    generate
    if ( USE_REG ) begin : ff_376
        reg   lut_376_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_376_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_376_ff <= lut_376_out;
            end
        end
        
        assign out_data[376] = lut_376_ff;
    end
    else begin : no_ff_376
        assign out_data[376] = lut_376_out;
    end
    endgenerate
    
    
    
    // LUT : 377
    wire [15:0] lut_377_table = 16'b1010101010101010;
    wire [3:0] lut_377_select = {
                             in_data[562],
                             in_data[71],
                             in_data[437],
                             in_data[313]};
    
    wire lut_377_out = lut_377_table[lut_377_select];
    
    generate
    if ( USE_REG ) begin : ff_377
        reg   lut_377_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_377_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_377_ff <= lut_377_out;
            end
        end
        
        assign out_data[377] = lut_377_ff;
    end
    else begin : no_ff_377
        assign out_data[377] = lut_377_out;
    end
    endgenerate
    
    
    
    // LUT : 378
    wire [15:0] lut_378_table = 16'b1111111111110101;
    wire [3:0] lut_378_select = {
                             in_data[618],
                             in_data[476],
                             in_data[91],
                             in_data[140]};
    
    wire lut_378_out = lut_378_table[lut_378_select];
    
    generate
    if ( USE_REG ) begin : ff_378
        reg   lut_378_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_378_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_378_ff <= lut_378_out;
            end
        end
        
        assign out_data[378] = lut_378_ff;
    end
    else begin : no_ff_378
        assign out_data[378] = lut_378_out;
    end
    endgenerate
    
    
    
    // LUT : 379
    wire [15:0] lut_379_table = 16'b1100111011000000;
    wire [3:0] lut_379_select = {
                             in_data[465],
                             in_data[251],
                             in_data[628],
                             in_data[322]};
    
    wire lut_379_out = lut_379_table[lut_379_select];
    
    generate
    if ( USE_REG ) begin : ff_379
        reg   lut_379_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_379_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_379_ff <= lut_379_out;
            end
        end
        
        assign out_data[379] = lut_379_ff;
    end
    else begin : no_ff_379
        assign out_data[379] = lut_379_out;
    end
    endgenerate
    
    
    
    // LUT : 380
    wire [15:0] lut_380_table = 16'b0010001010110011;
    wire [3:0] lut_380_select = {
                             in_data[625],
                             in_data[339],
                             in_data[452],
                             in_data[459]};
    
    wire lut_380_out = lut_380_table[lut_380_select];
    
    generate
    if ( USE_REG ) begin : ff_380
        reg   lut_380_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_380_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_380_ff <= lut_380_out;
            end
        end
        
        assign out_data[380] = lut_380_ff;
    end
    else begin : no_ff_380
        assign out_data[380] = lut_380_out;
    end
    endgenerate
    
    
    
    // LUT : 381
    wire [15:0] lut_381_table = 16'b1101110101001101;
    wire [3:0] lut_381_select = {
                             in_data[217],
                             in_data[455],
                             in_data[250],
                             in_data[14]};
    
    wire lut_381_out = lut_381_table[lut_381_select];
    
    generate
    if ( USE_REG ) begin : ff_381
        reg   lut_381_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_381_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_381_ff <= lut_381_out;
            end
        end
        
        assign out_data[381] = lut_381_ff;
    end
    else begin : no_ff_381
        assign out_data[381] = lut_381_out;
    end
    endgenerate
    
    
    
    // LUT : 382
    wire [15:0] lut_382_table = 16'b1000000011111111;
    wire [3:0] lut_382_select = {
                             in_data[359],
                             in_data[467],
                             in_data[67],
                             in_data[307]};
    
    wire lut_382_out = lut_382_table[lut_382_select];
    
    generate
    if ( USE_REG ) begin : ff_382
        reg   lut_382_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_382_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_382_ff <= lut_382_out;
            end
        end
        
        assign out_data[382] = lut_382_ff;
    end
    else begin : no_ff_382
        assign out_data[382] = lut_382_out;
    end
    endgenerate
    
    
    
    // LUT : 383
    wire [15:0] lut_383_table = 16'b1011001010111011;
    wire [3:0] lut_383_select = {
                             in_data[495],
                             in_data[109],
                             in_data[207],
                             in_data[555]};
    
    wire lut_383_out = lut_383_table[lut_383_select];
    
    generate
    if ( USE_REG ) begin : ff_383
        reg   lut_383_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_383_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_383_ff <= lut_383_out;
            end
        end
        
        assign out_data[383] = lut_383_ff;
    end
    else begin : no_ff_383
        assign out_data[383] = lut_383_out;
    end
    endgenerate
    
    
    
    // LUT : 384
    wire [15:0] lut_384_table = 16'b0101000001010101;
    wire [3:0] lut_384_select = {
                             in_data[297],
                             in_data[328],
                             in_data[360],
                             in_data[194]};
    
    wire lut_384_out = lut_384_table[lut_384_select];
    
    generate
    if ( USE_REG ) begin : ff_384
        reg   lut_384_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_384_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_384_ff <= lut_384_out;
            end
        end
        
        assign out_data[384] = lut_384_ff;
    end
    else begin : no_ff_384
        assign out_data[384] = lut_384_out;
    end
    endgenerate
    
    
    
    // LUT : 385
    wire [15:0] lut_385_table = 16'b0000001100110111;
    wire [3:0] lut_385_select = {
                             in_data[474],
                             in_data[24],
                             in_data[208],
                             in_data[128]};
    
    wire lut_385_out = lut_385_table[lut_385_select];
    
    generate
    if ( USE_REG ) begin : ff_385
        reg   lut_385_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_385_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_385_ff <= lut_385_out;
            end
        end
        
        assign out_data[385] = lut_385_ff;
    end
    else begin : no_ff_385
        assign out_data[385] = lut_385_out;
    end
    endgenerate
    
    
    
    // LUT : 386
    wire [15:0] lut_386_table = 16'b0011000111110001;
    wire [3:0] lut_386_select = {
                             in_data[257],
                             in_data[143],
                             in_data[382],
                             in_data[456]};
    
    wire lut_386_out = lut_386_table[lut_386_select];
    
    generate
    if ( USE_REG ) begin : ff_386
        reg   lut_386_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_386_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_386_ff <= lut_386_out;
            end
        end
        
        assign out_data[386] = lut_386_ff;
    end
    else begin : no_ff_386
        assign out_data[386] = lut_386_out;
    end
    endgenerate
    
    
    
    // LUT : 387
    wire [15:0] lut_387_table = 16'b0111010001000100;
    wire [3:0] lut_387_select = {
                             in_data[420],
                             in_data[185],
                             in_data[227],
                             in_data[617]};
    
    wire lut_387_out = lut_387_table[lut_387_select];
    
    generate
    if ( USE_REG ) begin : ff_387
        reg   lut_387_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_387_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_387_ff <= lut_387_out;
            end
        end
        
        assign out_data[387] = lut_387_ff;
    end
    else begin : no_ff_387
        assign out_data[387] = lut_387_out;
    end
    endgenerate
    
    
    
    // LUT : 388
    wire [15:0] lut_388_table = 16'b0000000010110011;
    wire [3:0] lut_388_select = {
                             in_data[177],
                             in_data[534],
                             in_data[285],
                             in_data[318]};
    
    wire lut_388_out = lut_388_table[lut_388_select];
    
    generate
    if ( USE_REG ) begin : ff_388
        reg   lut_388_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_388_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_388_ff <= lut_388_out;
            end
        end
        
        assign out_data[388] = lut_388_ff;
    end
    else begin : no_ff_388
        assign out_data[388] = lut_388_out;
    end
    endgenerate
    
    
    
    // LUT : 389
    wire [15:0] lut_389_table = 16'b0101111100000000;
    wire [3:0] lut_389_select = {
                             in_data[479],
                             in_data[175],
                             in_data[369],
                             in_data[54]};
    
    wire lut_389_out = lut_389_table[lut_389_select];
    
    generate
    if ( USE_REG ) begin : ff_389
        reg   lut_389_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_389_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_389_ff <= lut_389_out;
            end
        end
        
        assign out_data[389] = lut_389_ff;
    end
    else begin : no_ff_389
        assign out_data[389] = lut_389_out;
    end
    endgenerate
    
    
    
    // LUT : 390
    wire [15:0] lut_390_table = 16'b1100110101001100;
    wire [3:0] lut_390_select = {
                             in_data[43],
                             in_data[519],
                             in_data[388],
                             in_data[34]};
    
    wire lut_390_out = lut_390_table[lut_390_select];
    
    generate
    if ( USE_REG ) begin : ff_390
        reg   lut_390_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_390_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_390_ff <= lut_390_out;
            end
        end
        
        assign out_data[390] = lut_390_ff;
    end
    else begin : no_ff_390
        assign out_data[390] = lut_390_out;
    end
    endgenerate
    
    
    
    // LUT : 391
    wire [15:0] lut_391_table = 16'b1011000000000000;
    wire [3:0] lut_391_select = {
                             in_data[2],
                             in_data[301],
                             in_data[224],
                             in_data[567]};
    
    wire lut_391_out = lut_391_table[lut_391_select];
    
    generate
    if ( USE_REG ) begin : ff_391
        reg   lut_391_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_391_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_391_ff <= lut_391_out;
            end
        end
        
        assign out_data[391] = lut_391_ff;
    end
    else begin : no_ff_391
        assign out_data[391] = lut_391_out;
    end
    endgenerate
    
    
    
    // LUT : 392
    wire [15:0] lut_392_table = 16'b1111101010100000;
    wire [3:0] lut_392_select = {
                             in_data[440],
                             in_data[247],
                             in_data[220],
                             in_data[148]};
    
    wire lut_392_out = lut_392_table[lut_392_select];
    
    generate
    if ( USE_REG ) begin : ff_392
        reg   lut_392_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_392_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_392_ff <= lut_392_out;
            end
        end
        
        assign out_data[392] = lut_392_ff;
    end
    else begin : no_ff_392
        assign out_data[392] = lut_392_out;
    end
    endgenerate
    
    
    
    // LUT : 393
    wire [15:0] lut_393_table = 16'b1100000011101010;
    wire [3:0] lut_393_select = {
                             in_data[82],
                             in_data[117],
                             in_data[77],
                             in_data[179]};
    
    wire lut_393_out = lut_393_table[lut_393_select];
    
    generate
    if ( USE_REG ) begin : ff_393
        reg   lut_393_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_393_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_393_ff <= lut_393_out;
            end
        end
        
        assign out_data[393] = lut_393_ff;
    end
    else begin : no_ff_393
        assign out_data[393] = lut_393_out;
    end
    endgenerate
    
    
    
    // LUT : 394
    wire [15:0] lut_394_table = 16'b0000111100000111;
    wire [3:0] lut_394_select = {
                             in_data[264],
                             in_data[321],
                             in_data[46],
                             in_data[233]};
    
    wire lut_394_out = lut_394_table[lut_394_select];
    
    generate
    if ( USE_REG ) begin : ff_394
        reg   lut_394_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_394_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_394_ff <= lut_394_out;
            end
        end
        
        assign out_data[394] = lut_394_ff;
    end
    else begin : no_ff_394
        assign out_data[394] = lut_394_out;
    end
    endgenerate
    
    
    
    // LUT : 395
    wire [15:0] lut_395_table = 16'b1010101011111111;
    wire [3:0] lut_395_select = {
                             in_data[214],
                             in_data[12],
                             in_data[347],
                             in_data[103]};
    
    wire lut_395_out = lut_395_table[lut_395_select];
    
    generate
    if ( USE_REG ) begin : ff_395
        reg   lut_395_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_395_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_395_ff <= lut_395_out;
            end
        end
        
        assign out_data[395] = lut_395_ff;
    end
    else begin : no_ff_395
        assign out_data[395] = lut_395_out;
    end
    endgenerate
    
    
    
    // LUT : 396
    wire [15:0] lut_396_table = 16'b1100111100001111;
    wire [3:0] lut_396_select = {
                             in_data[244],
                             in_data[296],
                             in_data[497],
                             in_data[619]};
    
    wire lut_396_out = lut_396_table[lut_396_select];
    
    generate
    if ( USE_REG ) begin : ff_396
        reg   lut_396_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_396_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_396_ff <= lut_396_out;
            end
        end
        
        assign out_data[396] = lut_396_ff;
    end
    else begin : no_ff_396
        assign out_data[396] = lut_396_out;
    end
    endgenerate
    
    
    
    // LUT : 397
    wire [15:0] lut_397_table = 16'b1111110011101000;
    wire [3:0] lut_397_select = {
                             in_data[542],
                             in_data[606],
                             in_data[293],
                             in_data[520]};
    
    wire lut_397_out = lut_397_table[lut_397_select];
    
    generate
    if ( USE_REG ) begin : ff_397
        reg   lut_397_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_397_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_397_ff <= lut_397_out;
            end
        end
        
        assign out_data[397] = lut_397_ff;
    end
    else begin : no_ff_397
        assign out_data[397] = lut_397_out;
    end
    endgenerate
    
    
    
    // LUT : 398
    wire [15:0] lut_398_table = 16'b1111111100110000;
    wire [3:0] lut_398_select = {
                             in_data[575],
                             in_data[605],
                             in_data[65],
                             in_data[287]};
    
    wire lut_398_out = lut_398_table[lut_398_select];
    
    generate
    if ( USE_REG ) begin : ff_398
        reg   lut_398_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_398_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_398_ff <= lut_398_out;
            end
        end
        
        assign out_data[398] = lut_398_ff;
    end
    else begin : no_ff_398
        assign out_data[398] = lut_398_out;
    end
    endgenerate
    
    
    
    // LUT : 399
    wire [15:0] lut_399_table = 16'b0101111100000001;
    wire [3:0] lut_399_select = {
                             in_data[394],
                             in_data[601],
                             in_data[335],
                             in_data[445]};
    
    wire lut_399_out = lut_399_table[lut_399_select];
    
    generate
    if ( USE_REG ) begin : ff_399
        reg   lut_399_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_399_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_399_ff <= lut_399_out;
            end
        end
        
        assign out_data[399] = lut_399_ff;
    end
    else begin : no_ff_399
        assign out_data[399] = lut_399_out;
    end
    endgenerate
    
    
    
    // LUT : 400
    wire [15:0] lut_400_table = 16'b1110101011101010;
    wire [3:0] lut_400_select = {
                             in_data[237],
                             in_data[203],
                             in_data[212],
                             in_data[302]};
    
    wire lut_400_out = lut_400_table[lut_400_select];
    
    generate
    if ( USE_REG ) begin : ff_400
        reg   lut_400_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_400_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_400_ff <= lut_400_out;
            end
        end
        
        assign out_data[400] = lut_400_ff;
    end
    else begin : no_ff_400
        assign out_data[400] = lut_400_out;
    end
    endgenerate
    
    
    
    // LUT : 401
    wire [15:0] lut_401_table = 16'b0011101100000011;
    wire [3:0] lut_401_select = {
                             in_data[255],
                             in_data[88],
                             in_data[23],
                             in_data[422]};
    
    wire lut_401_out = lut_401_table[lut_401_select];
    
    generate
    if ( USE_REG ) begin : ff_401
        reg   lut_401_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_401_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_401_ff <= lut_401_out;
            end
        end
        
        assign out_data[401] = lut_401_ff;
    end
    else begin : no_ff_401
        assign out_data[401] = lut_401_out;
    end
    endgenerate
    
    
    
    // LUT : 402
    wire [15:0] lut_402_table = 16'b0011111100001111;
    wire [3:0] lut_402_select = {
                             in_data[401],
                             in_data[68],
                             in_data[7],
                             in_data[81]};
    
    wire lut_402_out = lut_402_table[lut_402_select];
    
    generate
    if ( USE_REG ) begin : ff_402
        reg   lut_402_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_402_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_402_ff <= lut_402_out;
            end
        end
        
        assign out_data[402] = lut_402_ff;
    end
    else begin : no_ff_402
        assign out_data[402] = lut_402_out;
    end
    endgenerate
    
    
    
    // LUT : 403
    wire [15:0] lut_403_table = 16'b0001111100000111;
    wire [3:0] lut_403_select = {
                             in_data[418],
                             in_data[95],
                             in_data[341],
                             in_data[130]};
    
    wire lut_403_out = lut_403_table[lut_403_select];
    
    generate
    if ( USE_REG ) begin : ff_403
        reg   lut_403_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_403_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_403_ff <= lut_403_out;
            end
        end
        
        assign out_data[403] = lut_403_ff;
    end
    else begin : no_ff_403
        assign out_data[403] = lut_403_out;
    end
    endgenerate
    
    
    
    // LUT : 404
    wire [15:0] lut_404_table = 16'b0001000100010001;
    wire [3:0] lut_404_select = {
                             in_data[271],
                             in_data[288],
                             in_data[19],
                             in_data[123]};
    
    wire lut_404_out = lut_404_table[lut_404_select];
    
    generate
    if ( USE_REG ) begin : ff_404
        reg   lut_404_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_404_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_404_ff <= lut_404_out;
            end
        end
        
        assign out_data[404] = lut_404_ff;
    end
    else begin : no_ff_404
        assign out_data[404] = lut_404_out;
    end
    endgenerate
    
    
    
    // LUT : 405
    wire [15:0] lut_405_table = 16'b1101111100000101;
    wire [3:0] lut_405_select = {
                             in_data[489],
                             in_data[131],
                             in_data[442],
                             in_data[549]};
    
    wire lut_405_out = lut_405_table[lut_405_select];
    
    generate
    if ( USE_REG ) begin : ff_405
        reg   lut_405_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_405_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_405_ff <= lut_405_out;
            end
        end
        
        assign out_data[405] = lut_405_ff;
    end
    else begin : no_ff_405
        assign out_data[405] = lut_405_out;
    end
    endgenerate
    
    
    
    // LUT : 406
    wire [15:0] lut_406_table = 16'b0111011101110111;
    wire [3:0] lut_406_select = {
                             in_data[229],
                             in_data[375],
                             in_data[379],
                             in_data[576]};
    
    wire lut_406_out = lut_406_table[lut_406_select];
    
    generate
    if ( USE_REG ) begin : ff_406
        reg   lut_406_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_406_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_406_ff <= lut_406_out;
            end
        end
        
        assign out_data[406] = lut_406_ff;
    end
    else begin : no_ff_406
        assign out_data[406] = lut_406_out;
    end
    endgenerate
    
    
    
    // LUT : 407
    wire [15:0] lut_407_table = 16'b0010001010101010;
    wire [3:0] lut_407_select = {
                             in_data[558],
                             in_data[323],
                             in_data[213],
                             in_data[20]};
    
    wire lut_407_out = lut_407_table[lut_407_select];
    
    generate
    if ( USE_REG ) begin : ff_407
        reg   lut_407_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_407_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_407_ff <= lut_407_out;
            end
        end
        
        assign out_data[407] = lut_407_ff;
    end
    else begin : no_ff_407
        assign out_data[407] = lut_407_out;
    end
    endgenerate
    
    
    
    // LUT : 408
    wire [15:0] lut_408_table = 16'b0011001101110011;
    wire [3:0] lut_408_select = {
                             in_data[9],
                             in_data[581],
                             in_data[320],
                             in_data[196]};
    
    wire lut_408_out = lut_408_table[lut_408_select];
    
    generate
    if ( USE_REG ) begin : ff_408
        reg   lut_408_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_408_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_408_ff <= lut_408_out;
            end
        end
        
        assign out_data[408] = lut_408_ff;
    end
    else begin : no_ff_408
        assign out_data[408] = lut_408_out;
    end
    endgenerate
    
    
    
    // LUT : 409
    wire [15:0] lut_409_table = 16'b0111001100110000;
    wire [3:0] lut_409_select = {
                             in_data[157],
                             in_data[566],
                             in_data[231],
                             in_data[309]};
    
    wire lut_409_out = lut_409_table[lut_409_select];
    
    generate
    if ( USE_REG ) begin : ff_409
        reg   lut_409_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_409_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_409_ff <= lut_409_out;
            end
        end
        
        assign out_data[409] = lut_409_ff;
    end
    else begin : no_ff_409
        assign out_data[409] = lut_409_out;
    end
    endgenerate
    
    
    
    // LUT : 410
    wire [15:0] lut_410_table = 16'b0011001100000010;
    wire [3:0] lut_410_select = {
                             in_data[319],
                             in_data[238],
                             in_data[28],
                             in_data[386]};
    
    wire lut_410_out = lut_410_table[lut_410_select];
    
    generate
    if ( USE_REG ) begin : ff_410
        reg   lut_410_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_410_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_410_ff <= lut_410_out;
            end
        end
        
        assign out_data[410] = lut_410_ff;
    end
    else begin : no_ff_410
        assign out_data[410] = lut_410_out;
    end
    endgenerate
    
    
    
    // LUT : 411
    wire [15:0] lut_411_table = 16'b1111000011110001;
    wire [3:0] lut_411_select = {
                             in_data[523],
                             in_data[639],
                             in_data[202],
                             in_data[331]};
    
    wire lut_411_out = lut_411_table[lut_411_select];
    
    generate
    if ( USE_REG ) begin : ff_411
        reg   lut_411_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_411_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_411_ff <= lut_411_out;
            end
        end
        
        assign out_data[411] = lut_411_ff;
    end
    else begin : no_ff_411
        assign out_data[411] = lut_411_out;
    end
    endgenerate
    
    
    
    // LUT : 412
    wire [15:0] lut_412_table = 16'b1101000001010000;
    wire [3:0] lut_412_select = {
                             in_data[522],
                             in_data[312],
                             in_data[350],
                             in_data[73]};
    
    wire lut_412_out = lut_412_table[lut_412_select];
    
    generate
    if ( USE_REG ) begin : ff_412
        reg   lut_412_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_412_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_412_ff <= lut_412_out;
            end
        end
        
        assign out_data[412] = lut_412_ff;
    end
    else begin : no_ff_412
        assign out_data[412] = lut_412_out;
    end
    endgenerate
    
    
    
    // LUT : 413
    wire [15:0] lut_413_table = 16'b0101010011010100;
    wire [3:0] lut_413_select = {
                             in_data[585],
                             in_data[326],
                             in_data[535],
                             in_data[571]};
    
    wire lut_413_out = lut_413_table[lut_413_select];
    
    generate
    if ( USE_REG ) begin : ff_413
        reg   lut_413_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_413_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_413_ff <= lut_413_out;
            end
        end
        
        assign out_data[413] = lut_413_ff;
    end
    else begin : no_ff_413
        assign out_data[413] = lut_413_out;
    end
    endgenerate
    
    
    
    // LUT : 414
    wire [15:0] lut_414_table = 16'b0111111100111111;
    wire [3:0] lut_414_select = {
                             in_data[594],
                             in_data[205],
                             in_data[514],
                             in_data[317]};
    
    wire lut_414_out = lut_414_table[lut_414_select];
    
    generate
    if ( USE_REG ) begin : ff_414
        reg   lut_414_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_414_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_414_ff <= lut_414_out;
            end
        end
        
        assign out_data[414] = lut_414_ff;
    end
    else begin : no_ff_414
        assign out_data[414] = lut_414_out;
    end
    endgenerate
    
    
    
    // LUT : 415
    wire [15:0] lut_415_table = 16'b0110110001110101;
    wire [3:0] lut_415_select = {
                             in_data[289],
                             in_data[547],
                             in_data[105],
                             in_data[589]};
    
    wire lut_415_out = lut_415_table[lut_415_select];
    
    generate
    if ( USE_REG ) begin : ff_415
        reg   lut_415_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_415_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_415_ff <= lut_415_out;
            end
        end
        
        assign out_data[415] = lut_415_ff;
    end
    else begin : no_ff_415
        assign out_data[415] = lut_415_out;
    end
    endgenerate
    
    
    
    // LUT : 416
    wire [15:0] lut_416_table = 16'b1010101011111011;
    wire [3:0] lut_416_select = {
                             in_data[416],
                             in_data[184],
                             in_data[115],
                             in_data[45]};
    
    wire lut_416_out = lut_416_table[lut_416_select];
    
    generate
    if ( USE_REG ) begin : ff_416
        reg   lut_416_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_416_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_416_ff <= lut_416_out;
            end
        end
        
        assign out_data[416] = lut_416_ff;
    end
    else begin : no_ff_416
        assign out_data[416] = lut_416_out;
    end
    endgenerate
    
    
    
    // LUT : 417
    wire [15:0] lut_417_table = 16'b1000100010001000;
    wire [3:0] lut_417_select = {
                             in_data[310],
                             in_data[76],
                             in_data[223],
                             in_data[336]};
    
    wire lut_417_out = lut_417_table[lut_417_select];
    
    generate
    if ( USE_REG ) begin : ff_417
        reg   lut_417_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_417_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_417_ff <= lut_417_out;
            end
        end
        
        assign out_data[417] = lut_417_ff;
    end
    else begin : no_ff_417
        assign out_data[417] = lut_417_out;
    end
    endgenerate
    
    
    
    // LUT : 418
    wire [15:0] lut_418_table = 16'b1111110011111000;
    wire [3:0] lut_418_select = {
                             in_data[259],
                             in_data[361],
                             in_data[15],
                             in_data[602]};
    
    wire lut_418_out = lut_418_table[lut_418_select];
    
    generate
    if ( USE_REG ) begin : ff_418
        reg   lut_418_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_418_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_418_ff <= lut_418_out;
            end
        end
        
        assign out_data[418] = lut_418_ff;
    end
    else begin : no_ff_418
        assign out_data[418] = lut_418_out;
    end
    endgenerate
    
    
    
    // LUT : 419
    wire [15:0] lut_419_table = 16'b0011001111111111;
    wire [3:0] lut_419_select = {
                             in_data[403],
                             in_data[475],
                             in_data[404],
                             in_data[92]};
    
    wire lut_419_out = lut_419_table[lut_419_select];
    
    generate
    if ( USE_REG ) begin : ff_419
        reg   lut_419_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_419_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_419_ff <= lut_419_out;
            end
        end
        
        assign out_data[419] = lut_419_ff;
    end
    else begin : no_ff_419
        assign out_data[419] = lut_419_out;
    end
    endgenerate
    
    
    
    // LUT : 420
    wire [15:0] lut_420_table = 16'b0011101100111011;
    wire [3:0] lut_420_select = {
                             in_data[596],
                             in_data[270],
                             in_data[161],
                             in_data[332]};
    
    wire lut_420_out = lut_420_table[lut_420_select];
    
    generate
    if ( USE_REG ) begin : ff_420
        reg   lut_420_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_420_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_420_ff <= lut_420_out;
            end
        end
        
        assign out_data[420] = lut_420_ff;
    end
    else begin : no_ff_420
        assign out_data[420] = lut_420_out;
    end
    endgenerate
    
    
    
    // LUT : 421
    wire [15:0] lut_421_table = 16'b0111001100110011;
    wire [3:0] lut_421_select = {
                             in_data[498],
                             in_data[541],
                             in_data[512],
                             in_data[572]};
    
    wire lut_421_out = lut_421_table[lut_421_select];
    
    generate
    if ( USE_REG ) begin : ff_421
        reg   lut_421_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_421_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_421_ff <= lut_421_out;
            end
        end
        
        assign out_data[421] = lut_421_ff;
    end
    else begin : no_ff_421
        assign out_data[421] = lut_421_out;
    end
    endgenerate
    
    
    
    // LUT : 422
    wire [15:0] lut_422_table = 16'b0011101100000000;
    wire [3:0] lut_422_select = {
                             in_data[254],
                             in_data[526],
                             in_data[84],
                             in_data[357]};
    
    wire lut_422_out = lut_422_table[lut_422_select];
    
    generate
    if ( USE_REG ) begin : ff_422
        reg   lut_422_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_422_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_422_ff <= lut_422_out;
            end
        end
        
        assign out_data[422] = lut_422_ff;
    end
    else begin : no_ff_422
        assign out_data[422] = lut_422_out;
    end
    endgenerate
    
    
    
    // LUT : 423
    wire [15:0] lut_423_table = 16'b1001101011111111;
    wire [3:0] lut_423_select = {
                             in_data[152],
                             in_data[482],
                             in_data[463],
                             in_data[574]};
    
    wire lut_423_out = lut_423_table[lut_423_select];
    
    generate
    if ( USE_REG ) begin : ff_423
        reg   lut_423_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_423_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_423_ff <= lut_423_out;
            end
        end
        
        assign out_data[423] = lut_423_ff;
    end
    else begin : no_ff_423
        assign out_data[423] = lut_423_out;
    end
    endgenerate
    
    
    
    // LUT : 424
    wire [15:0] lut_424_table = 16'b1111110111001101;
    wire [3:0] lut_424_select = {
                             in_data[496],
                             in_data[156],
                             in_data[169],
                             in_data[430]};
    
    wire lut_424_out = lut_424_table[lut_424_select];
    
    generate
    if ( USE_REG ) begin : ff_424
        reg   lut_424_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_424_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_424_ff <= lut_424_out;
            end
        end
        
        assign out_data[424] = lut_424_ff;
    end
    else begin : no_ff_424
        assign out_data[424] = lut_424_out;
    end
    endgenerate
    
    
    
    // LUT : 425
    wire [15:0] lut_425_table = 16'b1000100010000000;
    wire [3:0] lut_425_select = {
                             in_data[377],
                             in_data[348],
                             in_data[432],
                             in_data[218]};
    
    wire lut_425_out = lut_425_table[lut_425_select];
    
    generate
    if ( USE_REG ) begin : ff_425
        reg   lut_425_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_425_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_425_ff <= lut_425_out;
            end
        end
        
        assign out_data[425] = lut_425_ff;
    end
    else begin : no_ff_425
        assign out_data[425] = lut_425_out;
    end
    endgenerate
    
    
    
    // LUT : 426
    wire [15:0] lut_426_table = 16'b0000011100001011;
    wire [3:0] lut_426_select = {
                             in_data[537],
                             in_data[142],
                             in_data[358],
                             in_data[112]};
    
    wire lut_426_out = lut_426_table[lut_426_select];
    
    generate
    if ( USE_REG ) begin : ff_426
        reg   lut_426_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_426_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_426_ff <= lut_426_out;
            end
        end
        
        assign out_data[426] = lut_426_ff;
    end
    else begin : no_ff_426
        assign out_data[426] = lut_426_out;
    end
    endgenerate
    
    
    
    // LUT : 427
    wire [15:0] lut_427_table = 16'b1011111100000010;
    wire [3:0] lut_427_select = {
                             in_data[503],
                             in_data[485],
                             in_data[29],
                             in_data[536]};
    
    wire lut_427_out = lut_427_table[lut_427_select];
    
    generate
    if ( USE_REG ) begin : ff_427
        reg   lut_427_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_427_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_427_ff <= lut_427_out;
            end
        end
        
        assign out_data[427] = lut_427_ff;
    end
    else begin : no_ff_427
        assign out_data[427] = lut_427_out;
    end
    endgenerate
    
    
    
    // LUT : 428
    wire [15:0] lut_428_table = 16'b1011101100101010;
    wire [3:0] lut_428_select = {
                             in_data[508],
                             in_data[346],
                             in_data[491],
                             in_data[368]};
    
    wire lut_428_out = lut_428_table[lut_428_select];
    
    generate
    if ( USE_REG ) begin : ff_428
        reg   lut_428_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_428_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_428_ff <= lut_428_out;
            end
        end
        
        assign out_data[428] = lut_428_ff;
    end
    else begin : no_ff_428
        assign out_data[428] = lut_428_out;
    end
    endgenerate
    
    
    
    // LUT : 429
    wire [15:0] lut_429_table = 16'b1100000011001100;
    wire [3:0] lut_429_select = {
                             in_data[425],
                             in_data[191],
                             in_data[245],
                             in_data[144]};
    
    wire lut_429_out = lut_429_table[lut_429_select];
    
    generate
    if ( USE_REG ) begin : ff_429
        reg   lut_429_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_429_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_429_ff <= lut_429_out;
            end
        end
        
        assign out_data[429] = lut_429_ff;
    end
    else begin : no_ff_429
        assign out_data[429] = lut_429_out;
    end
    endgenerate
    
    
    
    // LUT : 430
    wire [15:0] lut_430_table = 16'b0000110101001100;
    wire [3:0] lut_430_select = {
                             in_data[620],
                             in_data[554],
                             in_data[515],
                             in_data[163]};
    
    wire lut_430_out = lut_430_table[lut_430_select];
    
    generate
    if ( USE_REG ) begin : ff_430
        reg   lut_430_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_430_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_430_ff <= lut_430_out;
            end
        end
        
        assign out_data[430] = lut_430_ff;
    end
    else begin : no_ff_430
        assign out_data[430] = lut_430_out;
    end
    endgenerate
    
    
    
    // LUT : 431
    wire [15:0] lut_431_table = 16'b0101100111111011;
    wire [3:0] lut_431_select = {
                             in_data[125],
                             in_data[635],
                             in_data[278],
                             in_data[395]};
    
    wire lut_431_out = lut_431_table[lut_431_select];
    
    generate
    if ( USE_REG ) begin : ff_431
        reg   lut_431_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_431_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_431_ff <= lut_431_out;
            end
        end
        
        assign out_data[431] = lut_431_ff;
    end
    else begin : no_ff_431
        assign out_data[431] = lut_431_out;
    end
    endgenerate
    
    
    
    // LUT : 432
    wire [15:0] lut_432_table = 16'b0100000101010111;
    wire [3:0] lut_432_select = {
                             in_data[171],
                             in_data[436],
                             in_data[390],
                             in_data[355]};
    
    wire lut_432_out = lut_432_table[lut_432_select];
    
    generate
    if ( USE_REG ) begin : ff_432
        reg   lut_432_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_432_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_432_ff <= lut_432_out;
            end
        end
        
        assign out_data[432] = lut_432_ff;
    end
    else begin : no_ff_432
        assign out_data[432] = lut_432_out;
    end
    endgenerate
    
    
    
    // LUT : 433
    wire [15:0] lut_433_table = 16'b1010000011111111;
    wire [3:0] lut_433_select = {
                             in_data[528],
                             in_data[444],
                             in_data[137],
                             in_data[316]};
    
    wire lut_433_out = lut_433_table[lut_433_select];
    
    generate
    if ( USE_REG ) begin : ff_433
        reg   lut_433_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_433_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_433_ff <= lut_433_out;
            end
        end
        
        assign out_data[433] = lut_433_ff;
    end
    else begin : no_ff_433
        assign out_data[433] = lut_433_out;
    end
    endgenerate
    
    
    
    // LUT : 434
    wire [15:0] lut_434_table = 16'b1111110111100000;
    wire [3:0] lut_434_select = {
                             in_data[372],
                             in_data[38],
                             in_data[187],
                             in_data[141]};
    
    wire lut_434_out = lut_434_table[lut_434_select];
    
    generate
    if ( USE_REG ) begin : ff_434
        reg   lut_434_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_434_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_434_ff <= lut_434_out;
            end
        end
        
        assign out_data[434] = lut_434_ff;
    end
    else begin : no_ff_434
        assign out_data[434] = lut_434_out;
    end
    endgenerate
    
    
    
    // LUT : 435
    wire [15:0] lut_435_table = 16'b1010100011101010;
    wire [3:0] lut_435_select = {
                             in_data[622],
                             in_data[85],
                             in_data[300],
                             in_data[234]};
    
    wire lut_435_out = lut_435_table[lut_435_select];
    
    generate
    if ( USE_REG ) begin : ff_435
        reg   lut_435_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_435_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_435_ff <= lut_435_out;
            end
        end
        
        assign out_data[435] = lut_435_ff;
    end
    else begin : no_ff_435
        assign out_data[435] = lut_435_out;
    end
    endgenerate
    
    
    
    // LUT : 436
    wire [15:0] lut_436_table = 16'b1010100010000000;
    wire [3:0] lut_436_select = {
                             in_data[344],
                             in_data[215],
                             in_data[488],
                             in_data[408]};
    
    wire lut_436_out = lut_436_table[lut_436_select];
    
    generate
    if ( USE_REG ) begin : ff_436
        reg   lut_436_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_436_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_436_ff <= lut_436_out;
            end
        end
        
        assign out_data[436] = lut_436_ff;
    end
    else begin : no_ff_436
        assign out_data[436] = lut_436_out;
    end
    endgenerate
    
    
    
    // LUT : 437
    wire [15:0] lut_437_table = 16'b1111000011110000;
    wire [3:0] lut_437_select = {
                             in_data[595],
                             in_data[94],
                             in_data[181],
                             in_data[461]};
    
    wire lut_437_out = lut_437_table[lut_437_select];
    
    generate
    if ( USE_REG ) begin : ff_437
        reg   lut_437_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_437_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_437_ff <= lut_437_out;
            end
        end
        
        assign out_data[437] = lut_437_ff;
    end
    else begin : no_ff_437
        assign out_data[437] = lut_437_out;
    end
    endgenerate
    
    
    
    // LUT : 438
    wire [15:0] lut_438_table = 16'b0101000111110111;
    wire [3:0] lut_438_select = {
                             in_data[120],
                             in_data[182],
                             in_data[334],
                             in_data[548]};
    
    wire lut_438_out = lut_438_table[lut_438_select];
    
    generate
    if ( USE_REG ) begin : ff_438
        reg   lut_438_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_438_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_438_ff <= lut_438_out;
            end
        end
        
        assign out_data[438] = lut_438_ff;
    end
    else begin : no_ff_438
        assign out_data[438] = lut_438_out;
    end
    endgenerate
    
    
    
    // LUT : 439
    wire [15:0] lut_439_table = 16'b0000010100000101;
    wire [3:0] lut_439_select = {
                             in_data[199],
                             in_data[4],
                             in_data[18],
                             in_data[183]};
    
    wire lut_439_out = lut_439_table[lut_439_select];
    
    generate
    if ( USE_REG ) begin : ff_439
        reg   lut_439_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_439_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_439_ff <= lut_439_out;
            end
        end
        
        assign out_data[439] = lut_439_ff;
    end
    else begin : no_ff_439
        assign out_data[439] = lut_439_out;
    end
    endgenerate
    
    
    
    // LUT : 440
    wire [15:0] lut_440_table = 16'b0010111100001011;
    wire [3:0] lut_440_select = {
                             in_data[158],
                             in_data[376],
                             in_data[116],
                             in_data[504]};
    
    wire lut_440_out = lut_440_table[lut_440_select];
    
    generate
    if ( USE_REG ) begin : ff_440
        reg   lut_440_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_440_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_440_ff <= lut_440_out;
            end
        end
        
        assign out_data[440] = lut_440_ff;
    end
    else begin : no_ff_440
        assign out_data[440] = lut_440_out;
    end
    endgenerate
    
    
    
    // LUT : 441
    wire [15:0] lut_441_table = 16'b0000000000100011;
    wire [3:0] lut_441_select = {
                             in_data[415],
                             in_data[417],
                             in_data[527],
                             in_data[494]};
    
    wire lut_441_out = lut_441_table[lut_441_select];
    
    generate
    if ( USE_REG ) begin : ff_441
        reg   lut_441_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_441_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_441_ff <= lut_441_out;
            end
        end
        
        assign out_data[441] = lut_441_ff;
    end
    else begin : no_ff_441
        assign out_data[441] = lut_441_out;
    end
    endgenerate
    
    
    
    // LUT : 442
    wire [15:0] lut_442_table = 16'b1101010101000000;
    wire [3:0] lut_442_select = {
                             in_data[530],
                             in_data[399],
                             in_data[352],
                             in_data[96]};
    
    wire lut_442_out = lut_442_table[lut_442_select];
    
    generate
    if ( USE_REG ) begin : ff_442
        reg   lut_442_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_442_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_442_ff <= lut_442_out;
            end
        end
        
        assign out_data[442] = lut_442_ff;
    end
    else begin : no_ff_442
        assign out_data[442] = lut_442_out;
    end
    endgenerate
    
    
    
    // LUT : 443
    wire [15:0] lut_443_table = 16'b1010101011101000;
    wire [3:0] lut_443_select = {
                             in_data[568],
                             in_data[275],
                             in_data[209],
                             in_data[127]};
    
    wire lut_443_out = lut_443_table[lut_443_select];
    
    generate
    if ( USE_REG ) begin : ff_443
        reg   lut_443_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_443_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_443_ff <= lut_443_out;
            end
        end
        
        assign out_data[443] = lut_443_ff;
    end
    else begin : no_ff_443
        assign out_data[443] = lut_443_out;
    end
    endgenerate
    
    
    
    // LUT : 444
    wire [15:0] lut_444_table = 16'b0010001000111011;
    wire [3:0] lut_444_select = {
                             in_data[57],
                             in_data[86],
                             in_data[343],
                             in_data[406]};
    
    wire lut_444_out = lut_444_table[lut_444_select];
    
    generate
    if ( USE_REG ) begin : ff_444
        reg   lut_444_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_444_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_444_ff <= lut_444_out;
            end
        end
        
        assign out_data[444] = lut_444_ff;
    end
    else begin : no_ff_444
        assign out_data[444] = lut_444_out;
    end
    endgenerate
    
    
    
    // LUT : 445
    wire [15:0] lut_445_table = 16'b1000101010101110;
    wire [3:0] lut_445_select = {
                             in_data[145],
                             in_data[64],
                             in_data[186],
                             in_data[22]};
    
    wire lut_445_out = lut_445_table[lut_445_select];
    
    generate
    if ( USE_REG ) begin : ff_445
        reg   lut_445_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_445_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_445_ff <= lut_445_out;
            end
        end
        
        assign out_data[445] = lut_445_ff;
    end
    else begin : no_ff_445
        assign out_data[445] = lut_445_out;
    end
    endgenerate
    
    
    
    // LUT : 446
    wire [15:0] lut_446_table = 16'b0111010100000000;
    wire [3:0] lut_446_select = {
                             in_data[201],
                             in_data[160],
                             in_data[546],
                             in_data[413]};
    
    wire lut_446_out = lut_446_table[lut_446_select];
    
    generate
    if ( USE_REG ) begin : ff_446
        reg   lut_446_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_446_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_446_ff <= lut_446_out;
            end
        end
        
        assign out_data[446] = lut_446_ff;
    end
    else begin : no_ff_446
        assign out_data[446] = lut_446_out;
    end
    endgenerate
    
    
    
    // LUT : 447
    wire [15:0] lut_447_table = 16'b1010000011111010;
    wire [3:0] lut_447_select = {
                             in_data[58],
                             in_data[383],
                             in_data[480],
                             in_data[342]};
    
    wire lut_447_out = lut_447_table[lut_447_select];
    
    generate
    if ( USE_REG ) begin : ff_447
        reg   lut_447_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_447_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_447_ff <= lut_447_out;
            end
        end
        
        assign out_data[447] = lut_447_ff;
    end
    else begin : no_ff_447
        assign out_data[447] = lut_447_out;
    end
    endgenerate
    
    
    
    // LUT : 448
    wire [15:0] lut_448_table = 16'b0001000101110011;
    wire [3:0] lut_448_select = {
                             in_data[41],
                             in_data[78],
                             in_data[545],
                             in_data[374]};
    
    wire lut_448_out = lut_448_table[lut_448_select];
    
    generate
    if ( USE_REG ) begin : ff_448
        reg   lut_448_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_448_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_448_ff <= lut_448_out;
            end
        end
        
        assign out_data[448] = lut_448_ff;
    end
    else begin : no_ff_448
        assign out_data[448] = lut_448_out;
    end
    endgenerate
    
    
    
    // LUT : 449
    wire [15:0] lut_449_table = 16'b0011001100100010;
    wire [3:0] lut_449_select = {
                             in_data[582],
                             in_data[172],
                             in_data[126],
                             in_data[102]};
    
    wire lut_449_out = lut_449_table[lut_449_select];
    
    generate
    if ( USE_REG ) begin : ff_449
        reg   lut_449_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_449_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_449_ff <= lut_449_out;
            end
        end
        
        assign out_data[449] = lut_449_ff;
    end
    else begin : no_ff_449
        assign out_data[449] = lut_449_out;
    end
    endgenerate
    
    
    
    // LUT : 450
    wire [15:0] lut_450_table = 16'b0001000100010001;
    wire [3:0] lut_450_select = {
                             in_data[99],
                             in_data[423],
                             in_data[32],
                             in_data[164]};
    
    wire lut_450_out = lut_450_table[lut_450_select];
    
    generate
    if ( USE_REG ) begin : ff_450
        reg   lut_450_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_450_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_450_ff <= lut_450_out;
            end
        end
        
        assign out_data[450] = lut_450_ff;
    end
    else begin : no_ff_450
        assign out_data[450] = lut_450_out;
    end
    endgenerate
    
    
    
    // LUT : 451
    wire [15:0] lut_451_table = 16'b0000000111011111;
    wire [3:0] lut_451_select = {
                             in_data[364],
                             in_data[139],
                             in_data[262],
                             in_data[265]};
    
    wire lut_451_out = lut_451_table[lut_451_select];
    
    generate
    if ( USE_REG ) begin : ff_451
        reg   lut_451_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_451_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_451_ff <= lut_451_out;
            end
        end
        
        assign out_data[451] = lut_451_ff;
    end
    else begin : no_ff_451
        assign out_data[451] = lut_451_out;
    end
    endgenerate
    
    
    
    // LUT : 452
    wire [15:0] lut_452_table = 16'b1100111010001110;
    wire [3:0] lut_452_select = {
                             in_data[613],
                             in_data[1],
                             in_data[155],
                             in_data[299]};
    
    wire lut_452_out = lut_452_table[lut_452_select];
    
    generate
    if ( USE_REG ) begin : ff_452
        reg   lut_452_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_452_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_452_ff <= lut_452_out;
            end
        end
        
        assign out_data[452] = lut_452_ff;
    end
    else begin : no_ff_452
        assign out_data[452] = lut_452_out;
    end
    endgenerate
    
    
    
    // LUT : 453
    wire [15:0] lut_453_table = 16'b1110111110001110;
    wire [3:0] lut_453_select = {
                             in_data[173],
                             in_data[10],
                             in_data[499],
                             in_data[69]};
    
    wire lut_453_out = lut_453_table[lut_453_select];
    
    generate
    if ( USE_REG ) begin : ff_453
        reg   lut_453_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_453_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_453_ff <= lut_453_out;
            end
        end
        
        assign out_data[453] = lut_453_ff;
    end
    else begin : no_ff_453
        assign out_data[453] = lut_453_out;
    end
    endgenerate
    
    
    
    // LUT : 454
    wire [15:0] lut_454_table = 16'b0010101010101111;
    wire [3:0] lut_454_select = {
                             in_data[431],
                             in_data[609],
                             in_data[384],
                             in_data[458]};
    
    wire lut_454_out = lut_454_table[lut_454_select];
    
    generate
    if ( USE_REG ) begin : ff_454
        reg   lut_454_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_454_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_454_ff <= lut_454_out;
            end
        end
        
        assign out_data[454] = lut_454_ff;
    end
    else begin : no_ff_454
        assign out_data[454] = lut_454_out;
    end
    endgenerate
    
    
    
    // LUT : 455
    wire [15:0] lut_455_table = 16'b1000101011111110;
    wire [3:0] lut_455_select = {
                             in_data[106],
                             in_data[48],
                             in_data[216],
                             in_data[441]};
    
    wire lut_455_out = lut_455_table[lut_455_select];
    
    generate
    if ( USE_REG ) begin : ff_455
        reg   lut_455_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_455_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_455_ff <= lut_455_out;
            end
        end
        
        assign out_data[455] = lut_455_ff;
    end
    else begin : no_ff_455
        assign out_data[455] = lut_455_out;
    end
    endgenerate
    
    
    
    // LUT : 456
    wire [15:0] lut_456_table = 16'b1100100011101111;
    wire [3:0] lut_456_select = {
                             in_data[240],
                             in_data[378],
                             in_data[427],
                             in_data[623]};
    
    wire lut_456_out = lut_456_table[lut_456_select];
    
    generate
    if ( USE_REG ) begin : ff_456
        reg   lut_456_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_456_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_456_ff <= lut_456_out;
            end
        end
        
        assign out_data[456] = lut_456_ff;
    end
    else begin : no_ff_456
        assign out_data[456] = lut_456_out;
    end
    endgenerate
    
    
    
    // LUT : 457
    wire [15:0] lut_457_table = 16'b1000100011111111;
    wire [3:0] lut_457_select = {
                             in_data[101],
                             in_data[314],
                             in_data[303],
                             in_data[435]};
    
    wire lut_457_out = lut_457_table[lut_457_select];
    
    generate
    if ( USE_REG ) begin : ff_457
        reg   lut_457_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_457_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_457_ff <= lut_457_out;
            end
        end
        
        assign out_data[457] = lut_457_ff;
    end
    else begin : no_ff_457
        assign out_data[457] = lut_457_out;
    end
    endgenerate
    
    
    
    // LUT : 458
    wire [15:0] lut_458_table = 16'b1100000011000000;
    wire [3:0] lut_458_select = {
                             in_data[393],
                             in_data[266],
                             in_data[189],
                             in_data[351]};
    
    wire lut_458_out = lut_458_table[lut_458_select];
    
    generate
    if ( USE_REG ) begin : ff_458
        reg   lut_458_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_458_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_458_ff <= lut_458_out;
            end
        end
        
        assign out_data[458] = lut_458_ff;
    end
    else begin : no_ff_458
        assign out_data[458] = lut_458_out;
    end
    endgenerate
    
    
    
    // LUT : 459
    wire [15:0] lut_459_table = 16'b0100000001011101;
    wire [3:0] lut_459_select = {
                             in_data[462],
                             in_data[228],
                             in_data[570],
                             in_data[63]};
    
    wire lut_459_out = lut_459_table[lut_459_select];
    
    generate
    if ( USE_REG ) begin : ff_459
        reg   lut_459_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_459_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_459_ff <= lut_459_out;
            end
        end
        
        assign out_data[459] = lut_459_ff;
    end
    else begin : no_ff_459
        assign out_data[459] = lut_459_out;
    end
    endgenerate
    
    
    
    // LUT : 460
    wire [15:0] lut_460_table = 16'b0000000011011111;
    wire [3:0] lut_460_select = {
                             in_data[614],
                             in_data[27],
                             in_data[354],
                             in_data[243]};
    
    wire lut_460_out = lut_460_table[lut_460_select];
    
    generate
    if ( USE_REG ) begin : ff_460
        reg   lut_460_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_460_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_460_ff <= lut_460_out;
            end
        end
        
        assign out_data[460] = lut_460_ff;
    end
    else begin : no_ff_460
        assign out_data[460] = lut_460_out;
    end
    endgenerate
    
    
    
    // LUT : 461
    wire [15:0] lut_461_table = 16'b1100110011101110;
    wire [3:0] lut_461_select = {
                             in_data[624],
                             in_data[525],
                             in_data[484],
                             in_data[89]};
    
    wire lut_461_out = lut_461_table[lut_461_select];
    
    generate
    if ( USE_REG ) begin : ff_461
        reg   lut_461_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_461_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_461_ff <= lut_461_out;
            end
        end
        
        assign out_data[461] = lut_461_ff;
    end
    else begin : no_ff_461
        assign out_data[461] = lut_461_out;
    end
    endgenerate
    
    
    
    // LUT : 462
    wire [15:0] lut_462_table = 16'b1100111111001111;
    wire [3:0] lut_462_select = {
                             in_data[481],
                             in_data[389],
                             in_data[146],
                             in_data[195]};
    
    wire lut_462_out = lut_462_table[lut_462_select];
    
    generate
    if ( USE_REG ) begin : ff_462
        reg   lut_462_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_462_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_462_ff <= lut_462_out;
            end
        end
        
        assign out_data[462] = lut_462_ff;
    end
    else begin : no_ff_462
        assign out_data[462] = lut_462_out;
    end
    endgenerate
    
    
    
    // LUT : 463
    wire [15:0] lut_463_table = 16'b1110111100000100;
    wire [3:0] lut_463_select = {
                             in_data[516],
                             in_data[42],
                             in_data[198],
                             in_data[210]};
    
    wire lut_463_out = lut_463_table[lut_463_select];
    
    generate
    if ( USE_REG ) begin : ff_463
        reg   lut_463_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_463_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_463_ff <= lut_463_out;
            end
        end
        
        assign out_data[463] = lut_463_ff;
    end
    else begin : no_ff_463
        assign out_data[463] = lut_463_out;
    end
    endgenerate
    
    
    
    // LUT : 464
    wire [15:0] lut_464_table = 16'b0011011100001111;
    wire [3:0] lut_464_select = {
                             in_data[402],
                             in_data[267],
                             in_data[236],
                             in_data[380]};
    
    wire lut_464_out = lut_464_table[lut_464_select];
    
    generate
    if ( USE_REG ) begin : ff_464
        reg   lut_464_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_464_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_464_ff <= lut_464_out;
            end
        end
        
        assign out_data[464] = lut_464_ff;
    end
    else begin : no_ff_464
        assign out_data[464] = lut_464_out;
    end
    endgenerate
    
    
    
    // LUT : 465
    wire [15:0] lut_465_table = 16'b0101010101010000;
    wire [3:0] lut_465_select = {
                             in_data[282],
                             in_data[483],
                             in_data[79],
                             in_data[363]};
    
    wire lut_465_out = lut_465_table[lut_465_select];
    
    generate
    if ( USE_REG ) begin : ff_465
        reg   lut_465_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_465_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_465_ff <= lut_465_out;
            end
        end
        
        assign out_data[465] = lut_465_ff;
    end
    else begin : no_ff_465
        assign out_data[465] = lut_465_out;
    end
    endgenerate
    
    
    
    // LUT : 466
    wire [15:0] lut_466_table = 16'b1101010111011101;
    wire [3:0] lut_466_select = {
                             in_data[249],
                             in_data[597],
                             in_data[340],
                             in_data[454]};
    
    wire lut_466_out = lut_466_table[lut_466_select];
    
    generate
    if ( USE_REG ) begin : ff_466
        reg   lut_466_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_466_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_466_ff <= lut_466_out;
            end
        end
        
        assign out_data[466] = lut_466_ff;
    end
    else begin : no_ff_466
        assign out_data[466] = lut_466_out;
    end
    endgenerate
    
    
    
    // LUT : 467
    wire [15:0] lut_467_table = 16'b1101110111000100;
    wire [3:0] lut_467_select = {
                             in_data[608],
                             in_data[226],
                             in_data[277],
                             in_data[241]};
    
    wire lut_467_out = lut_467_table[lut_467_select];
    
    generate
    if ( USE_REG ) begin : ff_467
        reg   lut_467_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_467_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_467_ff <= lut_467_out;
            end
        end
        
        assign out_data[467] = lut_467_ff;
    end
    else begin : no_ff_467
        assign out_data[467] = lut_467_out;
    end
    endgenerate
    
    
    
    // LUT : 468
    wire [15:0] lut_468_table = 16'b1000110011101110;
    wire [3:0] lut_468_select = {
                             in_data[100],
                             in_data[124],
                             in_data[400],
                             in_data[50]};
    
    wire lut_468_out = lut_468_table[lut_468_select];
    
    generate
    if ( USE_REG ) begin : ff_468
        reg   lut_468_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_468_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_468_ff <= lut_468_out;
            end
        end
        
        assign out_data[468] = lut_468_ff;
    end
    else begin : no_ff_468
        assign out_data[468] = lut_468_out;
    end
    endgenerate
    
    
    
    // LUT : 469
    wire [15:0] lut_469_table = 16'b0000110100001101;
    wire [3:0] lut_469_select = {
                             in_data[469],
                             in_data[17],
                             in_data[513],
                             in_data[118]};
    
    wire lut_469_out = lut_469_table[lut_469_select];
    
    generate
    if ( USE_REG ) begin : ff_469
        reg   lut_469_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_469_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_469_ff <= lut_469_out;
            end
        end
        
        assign out_data[469] = lut_469_ff;
    end
    else begin : no_ff_469
        assign out_data[469] = lut_469_out;
    end
    endgenerate
    
    
    
    // LUT : 470
    wire [15:0] lut_470_table = 16'b0000000100010011;
    wire [3:0] lut_470_select = {
                             in_data[630],
                             in_data[111],
                             in_data[66],
                             in_data[75]};
    
    wire lut_470_out = lut_470_table[lut_470_select];
    
    generate
    if ( USE_REG ) begin : ff_470
        reg   lut_470_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_470_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_470_ff <= lut_470_out;
            end
        end
        
        assign out_data[470] = lut_470_ff;
    end
    else begin : no_ff_470
        assign out_data[470] = lut_470_out;
    end
    endgenerate
    
    
    
    // LUT : 471
    wire [15:0] lut_471_table = 16'b0000101111111111;
    wire [3:0] lut_471_select = {
                             in_data[587],
                             in_data[439],
                             in_data[26],
                             in_data[391]};
    
    wire lut_471_out = lut_471_table[lut_471_select];
    
    generate
    if ( USE_REG ) begin : ff_471
        reg   lut_471_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_471_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_471_ff <= lut_471_out;
            end
        end
        
        assign out_data[471] = lut_471_ff;
    end
    else begin : no_ff_471
        assign out_data[471] = lut_471_out;
    end
    endgenerate
    
    
    
    // LUT : 472
    wire [15:0] lut_472_table = 16'b1111111100001000;
    wire [3:0] lut_472_select = {
                             in_data[239],
                             in_data[612],
                             in_data[3],
                             in_data[167]};
    
    wire lut_472_out = lut_472_table[lut_472_select];
    
    generate
    if ( USE_REG ) begin : ff_472
        reg   lut_472_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_472_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_472_ff <= lut_472_out;
            end
        end
        
        assign out_data[472] = lut_472_ff;
    end
    else begin : no_ff_472
        assign out_data[472] = lut_472_out;
    end
    endgenerate
    
    
    
    // LUT : 473
    wire [15:0] lut_473_table = 16'b0100000011011101;
    wire [3:0] lut_473_select = {
                             in_data[61],
                             in_data[412],
                             in_data[330],
                             in_data[252]};
    
    wire lut_473_out = lut_473_table[lut_473_select];
    
    generate
    if ( USE_REG ) begin : ff_473
        reg   lut_473_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_473_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_473_ff <= lut_473_out;
            end
        end
        
        assign out_data[473] = lut_473_ff;
    end
    else begin : no_ff_473
        assign out_data[473] = lut_473_out;
    end
    endgenerate
    
    
    
    // LUT : 474
    wire [15:0] lut_474_table = 16'b0000110011001100;
    wire [3:0] lut_474_select = {
                             in_data[563],
                             in_data[531],
                             in_data[586],
                             in_data[325]};
    
    wire lut_474_out = lut_474_table[lut_474_select];
    
    generate
    if ( USE_REG ) begin : ff_474
        reg   lut_474_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_474_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_474_ff <= lut_474_out;
            end
        end
        
        assign out_data[474] = lut_474_ff;
    end
    else begin : no_ff_474
        assign out_data[474] = lut_474_out;
    end
    endgenerate
    
    
    
    // LUT : 475
    wire [15:0] lut_475_table = 16'b0101110100001100;
    wire [3:0] lut_475_select = {
                             in_data[246],
                             in_data[135],
                             in_data[472],
                             in_data[33]};
    
    wire lut_475_out = lut_475_table[lut_475_select];
    
    generate
    if ( USE_REG ) begin : ff_475
        reg   lut_475_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_475_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_475_ff <= lut_475_out;
            end
        end
        
        assign out_data[475] = lut_475_ff;
    end
    else begin : no_ff_475
        assign out_data[475] = lut_475_out;
    end
    endgenerate
    
    
    
    // LUT : 476
    wire [15:0] lut_476_table = 16'b0101011100000011;
    wire [3:0] lut_476_select = {
                             in_data[221],
                             in_data[87],
                             in_data[371],
                             in_data[577]};
    
    wire lut_476_out = lut_476_table[lut_476_select];
    
    generate
    if ( USE_REG ) begin : ff_476
        reg   lut_476_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_476_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_476_ff <= lut_476_out;
            end
        end
        
        assign out_data[476] = lut_476_ff;
    end
    else begin : no_ff_476
        assign out_data[476] = lut_476_out;
    end
    endgenerate
    
    
    
    // LUT : 477
    wire [15:0] lut_477_table = 16'b0000100000001111;
    wire [3:0] lut_477_select = {
                             in_data[510],
                             in_data[457],
                             in_data[598],
                             in_data[593]};
    
    wire lut_477_out = lut_477_table[lut_477_select];
    
    generate
    if ( USE_REG ) begin : ff_477
        reg   lut_477_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_477_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_477_ff <= lut_477_out;
            end
        end
        
        assign out_data[477] = lut_477_ff;
    end
    else begin : no_ff_477
        assign out_data[477] = lut_477_out;
    end
    endgenerate
    
    
    
    // LUT : 478
    wire [15:0] lut_478_table = 16'b0010101010111111;
    wire [3:0] lut_478_select = {
                             in_data[592],
                             in_data[373],
                             in_data[551],
                             in_data[543]};
    
    wire lut_478_out = lut_478_table[lut_478_select];
    
    generate
    if ( USE_REG ) begin : ff_478
        reg   lut_478_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_478_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_478_ff <= lut_478_out;
            end
        end
        
        assign out_data[478] = lut_478_ff;
    end
    else begin : no_ff_478
        assign out_data[478] = lut_478_out;
    end
    endgenerate
    
    
    
    // LUT : 479
    wire [15:0] lut_479_table = 16'b1010101110101010;
    wire [3:0] lut_479_select = {
                             in_data[532],
                             in_data[72],
                             in_data[269],
                             in_data[178]};
    
    wire lut_479_out = lut_479_table[lut_479_select];
    
    generate
    if ( USE_REG ) begin : ff_479
        reg   lut_479_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_479_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_479_ff <= lut_479_out;
            end
        end
        
        assign out_data[479] = lut_479_ff;
    end
    else begin : no_ff_479
        assign out_data[479] = lut_479_out;
    end
    endgenerate
    
    
    
    // LUT : 480
    wire [15:0] lut_480_table = 16'b0000111100011111;
    wire [3:0] lut_480_select = {
                             in_data[103],
                             in_data[294],
                             in_data[634],
                             in_data[472]};
    
    wire lut_480_out = lut_480_table[lut_480_select];
    
    generate
    if ( USE_REG ) begin : ff_480
        reg   lut_480_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_480_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_480_ff <= lut_480_out;
            end
        end
        
        assign out_data[480] = lut_480_ff;
    end
    else begin : no_ff_480
        assign out_data[480] = lut_480_out;
    end
    endgenerate
    
    
    
    // LUT : 481
    wire [15:0] lut_481_table = 16'b1111101100110011;
    wire [3:0] lut_481_select = {
                             in_data[68],
                             in_data[444],
                             in_data[513],
                             in_data[332]};
    
    wire lut_481_out = lut_481_table[lut_481_select];
    
    generate
    if ( USE_REG ) begin : ff_481
        reg   lut_481_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_481_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_481_ff <= lut_481_out;
            end
        end
        
        assign out_data[481] = lut_481_ff;
    end
    else begin : no_ff_481
        assign out_data[481] = lut_481_out;
    end
    endgenerate
    
    
    
    // LUT : 482
    wire [15:0] lut_482_table = 16'b0101010111011111;
    wire [3:0] lut_482_select = {
                             in_data[461],
                             in_data[46],
                             in_data[35],
                             in_data[88]};
    
    wire lut_482_out = lut_482_table[lut_482_select];
    
    generate
    if ( USE_REG ) begin : ff_482
        reg   lut_482_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_482_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_482_ff <= lut_482_out;
            end
        end
        
        assign out_data[482] = lut_482_ff;
    end
    else begin : no_ff_482
        assign out_data[482] = lut_482_out;
    end
    endgenerate
    
    
    
    // LUT : 483
    wire [15:0] lut_483_table = 16'b1100000011000100;
    wire [3:0] lut_483_select = {
                             in_data[143],
                             in_data[504],
                             in_data[375],
                             in_data[39]};
    
    wire lut_483_out = lut_483_table[lut_483_select];
    
    generate
    if ( USE_REG ) begin : ff_483
        reg   lut_483_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_483_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_483_ff <= lut_483_out;
            end
        end
        
        assign out_data[483] = lut_483_ff;
    end
    else begin : no_ff_483
        assign out_data[483] = lut_483_out;
    end
    endgenerate
    
    
    
    // LUT : 484
    wire [15:0] lut_484_table = 16'b1111111100001111;
    wire [3:0] lut_484_select = {
                             in_data[267],
                             in_data[601],
                             in_data[628],
                             in_data[414]};
    
    wire lut_484_out = lut_484_table[lut_484_select];
    
    generate
    if ( USE_REG ) begin : ff_484
        reg   lut_484_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_484_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_484_ff <= lut_484_out;
            end
        end
        
        assign out_data[484] = lut_484_ff;
    end
    else begin : no_ff_484
        assign out_data[484] = lut_484_out;
    end
    endgenerate
    
    
    
    // LUT : 485
    wire [15:0] lut_485_table = 16'b0111011100110001;
    wire [3:0] lut_485_select = {
                             in_data[142],
                             in_data[200],
                             in_data[521],
                             in_data[223]};
    
    wire lut_485_out = lut_485_table[lut_485_select];
    
    generate
    if ( USE_REG ) begin : ff_485
        reg   lut_485_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_485_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_485_ff <= lut_485_out;
            end
        end
        
        assign out_data[485] = lut_485_ff;
    end
    else begin : no_ff_485
        assign out_data[485] = lut_485_out;
    end
    endgenerate
    
    
    
    // LUT : 486
    wire [15:0] lut_486_table = 16'b1111010111110101;
    wire [3:0] lut_486_select = {
                             in_data[542],
                             in_data[44],
                             in_data[333],
                             in_data[576]};
    
    wire lut_486_out = lut_486_table[lut_486_select];
    
    generate
    if ( USE_REG ) begin : ff_486
        reg   lut_486_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_486_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_486_ff <= lut_486_out;
            end
        end
        
        assign out_data[486] = lut_486_ff;
    end
    else begin : no_ff_486
        assign out_data[486] = lut_486_out;
    end
    endgenerate
    
    
    
    // LUT : 487
    wire [15:0] lut_487_table = 16'b1111111111001000;
    wire [3:0] lut_487_select = {
                             in_data[41],
                             in_data[522],
                             in_data[290],
                             in_data[323]};
    
    wire lut_487_out = lut_487_table[lut_487_select];
    
    generate
    if ( USE_REG ) begin : ff_487
        reg   lut_487_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_487_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_487_ff <= lut_487_out;
            end
        end
        
        assign out_data[487] = lut_487_ff;
    end
    else begin : no_ff_487
        assign out_data[487] = lut_487_out;
    end
    endgenerate
    
    
    
    // LUT : 488
    wire [15:0] lut_488_table = 16'b1010101000000000;
    wire [3:0] lut_488_select = {
                             in_data[297],
                             in_data[2],
                             in_data[562],
                             in_data[626]};
    
    wire lut_488_out = lut_488_table[lut_488_select];
    
    generate
    if ( USE_REG ) begin : ff_488
        reg   lut_488_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_488_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_488_ff <= lut_488_out;
            end
        end
        
        assign out_data[488] = lut_488_ff;
    end
    else begin : no_ff_488
        assign out_data[488] = lut_488_out;
    end
    endgenerate
    
    
    
    // LUT : 489
    wire [15:0] lut_489_table = 16'b1000110010001100;
    wire [3:0] lut_489_select = {
                             in_data[558],
                             in_data[228],
                             in_data[439],
                             in_data[572]};
    
    wire lut_489_out = lut_489_table[lut_489_select];
    
    generate
    if ( USE_REG ) begin : ff_489
        reg   lut_489_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_489_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_489_ff <= lut_489_out;
            end
        end
        
        assign out_data[489] = lut_489_ff;
    end
    else begin : no_ff_489
        assign out_data[489] = lut_489_out;
    end
    endgenerate
    
    
    
    // LUT : 490
    wire [15:0] lut_490_table = 16'b0011000011111111;
    wire [3:0] lut_490_select = {
                             in_data[420],
                             in_data[28],
                             in_data[604],
                             in_data[78]};
    
    wire lut_490_out = lut_490_table[lut_490_select];
    
    generate
    if ( USE_REG ) begin : ff_490
        reg   lut_490_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_490_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_490_ff <= lut_490_out;
            end
        end
        
        assign out_data[490] = lut_490_ff;
    end
    else begin : no_ff_490
        assign out_data[490] = lut_490_out;
    end
    endgenerate
    
    
    
    // LUT : 491
    wire [15:0] lut_491_table = 16'b0001000001110000;
    wire [3:0] lut_491_select = {
                             in_data[496],
                             in_data[274],
                             in_data[411],
                             in_data[520]};
    
    wire lut_491_out = lut_491_table[lut_491_select];
    
    generate
    if ( USE_REG ) begin : ff_491
        reg   lut_491_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_491_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_491_ff <= lut_491_out;
            end
        end
        
        assign out_data[491] = lut_491_ff;
    end
    else begin : no_ff_491
        assign out_data[491] = lut_491_out;
    end
    endgenerate
    
    
    
    // LUT : 492
    wire [15:0] lut_492_table = 16'b1100111111001111;
    wire [3:0] lut_492_select = {
                             in_data[292],
                             in_data[112],
                             in_data[340],
                             in_data[557]};
    
    wire lut_492_out = lut_492_table[lut_492_select];
    
    generate
    if ( USE_REG ) begin : ff_492
        reg   lut_492_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_492_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_492_ff <= lut_492_out;
            end
        end
        
        assign out_data[492] = lut_492_ff;
    end
    else begin : no_ff_492
        assign out_data[492] = lut_492_out;
    end
    endgenerate
    
    
    
    // LUT : 493
    wire [15:0] lut_493_table = 16'b0101010100000100;
    wire [3:0] lut_493_select = {
                             in_data[239],
                             in_data[402],
                             in_data[624],
                             in_data[61]};
    
    wire lut_493_out = lut_493_table[lut_493_select];
    
    generate
    if ( USE_REG ) begin : ff_493
        reg   lut_493_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_493_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_493_ff <= lut_493_out;
            end
        end
        
        assign out_data[493] = lut_493_ff;
    end
    else begin : no_ff_493
        assign out_data[493] = lut_493_out;
    end
    endgenerate
    
    
    
    // LUT : 494
    wire [15:0] lut_494_table = 16'b1110111011101110;
    wire [3:0] lut_494_select = {
                             in_data[413],
                             in_data[567],
                             in_data[91],
                             in_data[426]};
    
    wire lut_494_out = lut_494_table[lut_494_select];
    
    generate
    if ( USE_REG ) begin : ff_494
        reg   lut_494_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_494_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_494_ff <= lut_494_out;
            end
        end
        
        assign out_data[494] = lut_494_ff;
    end
    else begin : no_ff_494
        assign out_data[494] = lut_494_out;
    end
    endgenerate
    
    
    
    // LUT : 495
    wire [15:0] lut_495_table = 16'b0011000111110011;
    wire [3:0] lut_495_select = {
                             in_data[531],
                             in_data[174],
                             in_data[328],
                             in_data[638]};
    
    wire lut_495_out = lut_495_table[lut_495_select];
    
    generate
    if ( USE_REG ) begin : ff_495
        reg   lut_495_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_495_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_495_ff <= lut_495_out;
            end
        end
        
        assign out_data[495] = lut_495_ff;
    end
    else begin : no_ff_495
        assign out_data[495] = lut_495_out;
    end
    endgenerate
    
    
    
    // LUT : 496
    wire [15:0] lut_496_table = 16'b0101111100001111;
    wire [3:0] lut_496_select = {
                             in_data[145],
                             in_data[101],
                             in_data[373],
                             in_data[410]};
    
    wire lut_496_out = lut_496_table[lut_496_select];
    
    generate
    if ( USE_REG ) begin : ff_496
        reg   lut_496_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_496_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_496_ff <= lut_496_out;
            end
        end
        
        assign out_data[496] = lut_496_ff;
    end
    else begin : no_ff_496
        assign out_data[496] = lut_496_out;
    end
    endgenerate
    
    
    
    // LUT : 497
    wire [15:0] lut_497_table = 16'b1111011000100000;
    wire [3:0] lut_497_select = {
                             in_data[178],
                             in_data[617],
                             in_data[519],
                             in_data[453]};
    
    wire lut_497_out = lut_497_table[lut_497_select];
    
    generate
    if ( USE_REG ) begin : ff_497
        reg   lut_497_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_497_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_497_ff <= lut_497_out;
            end
        end
        
        assign out_data[497] = lut_497_ff;
    end
    else begin : no_ff_497
        assign out_data[497] = lut_497_out;
    end
    endgenerate
    
    
    
    // LUT : 498
    wire [15:0] lut_498_table = 16'b1010000010111011;
    wire [3:0] lut_498_select = {
                             in_data[72],
                             in_data[552],
                             in_data[443],
                             in_data[246]};
    
    wire lut_498_out = lut_498_table[lut_498_select];
    
    generate
    if ( USE_REG ) begin : ff_498
        reg   lut_498_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_498_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_498_ff <= lut_498_out;
            end
        end
        
        assign out_data[498] = lut_498_ff;
    end
    else begin : no_ff_498
        assign out_data[498] = lut_498_out;
    end
    endgenerate
    
    
    
    // LUT : 499
    wire [15:0] lut_499_table = 16'b1010101000001000;
    wire [3:0] lut_499_select = {
                             in_data[425],
                             in_data[462],
                             in_data[157],
                             in_data[586]};
    
    wire lut_499_out = lut_499_table[lut_499_select];
    
    generate
    if ( USE_REG ) begin : ff_499
        reg   lut_499_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_499_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_499_ff <= lut_499_out;
            end
        end
        
        assign out_data[499] = lut_499_ff;
    end
    else begin : no_ff_499
        assign out_data[499] = lut_499_out;
    end
    endgenerate
    
    
    
    // LUT : 500
    wire [15:0] lut_500_table = 16'b0111001100110000;
    wire [3:0] lut_500_select = {
                             in_data[129],
                             in_data[465],
                             in_data[484],
                             in_data[170]};
    
    wire lut_500_out = lut_500_table[lut_500_select];
    
    generate
    if ( USE_REG ) begin : ff_500
        reg   lut_500_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_500_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_500_ff <= lut_500_out;
            end
        end
        
        assign out_data[500] = lut_500_ff;
    end
    else begin : no_ff_500
        assign out_data[500] = lut_500_out;
    end
    endgenerate
    
    
    
    // LUT : 501
    wire [15:0] lut_501_table = 16'b0111011101010001;
    wire [3:0] lut_501_select = {
                             in_data[321],
                             in_data[59],
                             in_data[302],
                             in_data[264]};
    
    wire lut_501_out = lut_501_table[lut_501_select];
    
    generate
    if ( USE_REG ) begin : ff_501
        reg   lut_501_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_501_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_501_ff <= lut_501_out;
            end
        end
        
        assign out_data[501] = lut_501_ff;
    end
    else begin : no_ff_501
        assign out_data[501] = lut_501_out;
    end
    endgenerate
    
    
    
    // LUT : 502
    wire [15:0] lut_502_table = 16'b0101111100000001;
    wire [3:0] lut_502_select = {
                             in_data[283],
                             in_data[349],
                             in_data[573],
                             in_data[564]};
    
    wire lut_502_out = lut_502_table[lut_502_select];
    
    generate
    if ( USE_REG ) begin : ff_502
        reg   lut_502_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_502_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_502_ff <= lut_502_out;
            end
        end
        
        assign out_data[502] = lut_502_ff;
    end
    else begin : no_ff_502
        assign out_data[502] = lut_502_out;
    end
    endgenerate
    
    
    
    // LUT : 503
    wire [15:0] lut_503_table = 16'b1100110111000100;
    wire [3:0] lut_503_select = {
                             in_data[151],
                             in_data[6],
                             in_data[155],
                             in_data[140]};
    
    wire lut_503_out = lut_503_table[lut_503_select];
    
    generate
    if ( USE_REG ) begin : ff_503
        reg   lut_503_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_503_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_503_ff <= lut_503_out;
            end
        end
        
        assign out_data[503] = lut_503_ff;
    end
    else begin : no_ff_503
        assign out_data[503] = lut_503_out;
    end
    endgenerate
    
    
    
    // LUT : 504
    wire [15:0] lut_504_table = 16'b0001000101010001;
    wire [3:0] lut_504_select = {
                             in_data[296],
                             in_data[540],
                             in_data[547],
                             in_data[251]};
    
    wire lut_504_out = lut_504_table[lut_504_select];
    
    generate
    if ( USE_REG ) begin : ff_504
        reg   lut_504_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_504_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_504_ff <= lut_504_out;
            end
        end
        
        assign out_data[504] = lut_504_ff;
    end
    else begin : no_ff_504
        assign out_data[504] = lut_504_out;
    end
    endgenerate
    
    
    
    // LUT : 505
    wire [15:0] lut_505_table = 16'b1110111110001010;
    wire [3:0] lut_505_select = {
                             in_data[190],
                             in_data[185],
                             in_data[368],
                             in_data[516]};
    
    wire lut_505_out = lut_505_table[lut_505_select];
    
    generate
    if ( USE_REG ) begin : ff_505
        reg   lut_505_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_505_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_505_ff <= lut_505_out;
            end
        end
        
        assign out_data[505] = lut_505_ff;
    end
    else begin : no_ff_505
        assign out_data[505] = lut_505_out;
    end
    endgenerate
    
    
    
    // LUT : 506
    wire [15:0] lut_506_table = 16'b0011111100010000;
    wire [3:0] lut_506_select = {
                             in_data[153],
                             in_data[478],
                             in_data[172],
                             in_data[199]};
    
    wire lut_506_out = lut_506_table[lut_506_select];
    
    generate
    if ( USE_REG ) begin : ff_506
        reg   lut_506_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_506_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_506_ff <= lut_506_out;
            end
        end
        
        assign out_data[506] = lut_506_ff;
    end
    else begin : no_ff_506
        assign out_data[506] = lut_506_out;
    end
    endgenerate
    
    
    
    // LUT : 507
    wire [15:0] lut_507_table = 16'b1101010011000000;
    wire [3:0] lut_507_select = {
                             in_data[236],
                             in_data[389],
                             in_data[249],
                             in_data[227]};
    
    wire lut_507_out = lut_507_table[lut_507_select];
    
    generate
    if ( USE_REG ) begin : ff_507
        reg   lut_507_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_507_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_507_ff <= lut_507_out;
            end
        end
        
        assign out_data[507] = lut_507_ff;
    end
    else begin : no_ff_507
        assign out_data[507] = lut_507_out;
    end
    endgenerate
    
    
    
    // LUT : 508
    wire [15:0] lut_508_table = 16'b0001000100110111;
    wire [3:0] lut_508_select = {
                             in_data[127],
                             in_data[130],
                             in_data[337],
                             in_data[10]};
    
    wire lut_508_out = lut_508_table[lut_508_select];
    
    generate
    if ( USE_REG ) begin : ff_508
        reg   lut_508_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_508_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_508_ff <= lut_508_out;
            end
        end
        
        assign out_data[508] = lut_508_ff;
    end
    else begin : no_ff_508
        assign out_data[508] = lut_508_out;
    end
    endgenerate
    
    
    
    // LUT : 509
    wire [15:0] lut_509_table = 16'b1111000011111111;
    wire [3:0] lut_509_select = {
                             in_data[204],
                             in_data[416],
                             in_data[448],
                             in_data[639]};
    
    wire lut_509_out = lut_509_table[lut_509_select];
    
    generate
    if ( USE_REG ) begin : ff_509
        reg   lut_509_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_509_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_509_ff <= lut_509_out;
            end
        end
        
        assign out_data[509] = lut_509_ff;
    end
    else begin : no_ff_509
        assign out_data[509] = lut_509_out;
    end
    endgenerate
    
    
    
    // LUT : 510
    wire [15:0] lut_510_table = 16'b0000111100000111;
    wire [3:0] lut_510_select = {
                             in_data[355],
                             in_data[511],
                             in_data[554],
                             in_data[445]};
    
    wire lut_510_out = lut_510_table[lut_510_select];
    
    generate
    if ( USE_REG ) begin : ff_510
        reg   lut_510_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_510_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_510_ff <= lut_510_out;
            end
        end
        
        assign out_data[510] = lut_510_ff;
    end
    else begin : no_ff_510
        assign out_data[510] = lut_510_out;
    end
    endgenerate
    
    
    
    // LUT : 511
    wire [15:0] lut_511_table = 16'b0010001010111011;
    wire [3:0] lut_511_select = {
                             in_data[360],
                             in_data[109],
                             in_data[419],
                             in_data[0]};
    
    wire lut_511_out = lut_511_table[lut_511_select];
    
    generate
    if ( USE_REG ) begin : ff_511
        reg   lut_511_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_511_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_511_ff <= lut_511_out;
            end
        end
        
        assign out_data[511] = lut_511_ff;
    end
    else begin : no_ff_511
        assign out_data[511] = lut_511_out;
    end
    endgenerate
    
    
    
    // LUT : 512
    wire [15:0] lut_512_table = 16'b0001000011110101;
    wire [3:0] lut_512_select = {
                             in_data[73],
                             in_data[134],
                             in_data[481],
                             in_data[235]};
    
    wire lut_512_out = lut_512_table[lut_512_select];
    
    generate
    if ( USE_REG ) begin : ff_512
        reg   lut_512_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_512_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_512_ff <= lut_512_out;
            end
        end
        
        assign out_data[512] = lut_512_ff;
    end
    else begin : no_ff_512
        assign out_data[512] = lut_512_out;
    end
    endgenerate
    
    
    
    // LUT : 513
    wire [15:0] lut_513_table = 16'b0010001000100010;
    wire [3:0] lut_513_select = {
                             in_data[180],
                             in_data[238],
                             in_data[596],
                             in_data[5]};
    
    wire lut_513_out = lut_513_table[lut_513_select];
    
    generate
    if ( USE_REG ) begin : ff_513
        reg   lut_513_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_513_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_513_ff <= lut_513_out;
            end
        end
        
        assign out_data[513] = lut_513_ff;
    end
    else begin : no_ff_513
        assign out_data[513] = lut_513_out;
    end
    endgenerate
    
    
    
    // LUT : 514
    wire [15:0] lut_514_table = 16'b0000000011101100;
    wire [3:0] lut_514_select = {
                             in_data[629],
                             in_data[125],
                             in_data[428],
                             in_data[591]};
    
    wire lut_514_out = lut_514_table[lut_514_select];
    
    generate
    if ( USE_REG ) begin : ff_514
        reg   lut_514_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_514_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_514_ff <= lut_514_out;
            end
        end
        
        assign out_data[514] = lut_514_ff;
    end
    else begin : no_ff_514
        assign out_data[514] = lut_514_out;
    end
    endgenerate
    
    
    
    // LUT : 515
    wire [15:0] lut_515_table = 16'b0001000011110011;
    wire [3:0] lut_515_select = {
                             in_data[133],
                             in_data[118],
                             in_data[14],
                             in_data[255]};
    
    wire lut_515_out = lut_515_table[lut_515_select];
    
    generate
    if ( USE_REG ) begin : ff_515
        reg   lut_515_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_515_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_515_ff <= lut_515_out;
            end
        end
        
        assign out_data[515] = lut_515_ff;
    end
    else begin : no_ff_515
        assign out_data[515] = lut_515_out;
    end
    endgenerate
    
    
    
    // LUT : 516
    wire [15:0] lut_516_table = 16'b0100100000001110;
    wire [3:0] lut_516_select = {
                             in_data[363],
                             in_data[148],
                             in_data[300],
                             in_data[268]};
    
    wire lut_516_out = lut_516_table[lut_516_select];
    
    generate
    if ( USE_REG ) begin : ff_516
        reg   lut_516_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_516_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_516_ff <= lut_516_out;
            end
        end
        
        assign out_data[516] = lut_516_ff;
    end
    else begin : no_ff_516
        assign out_data[516] = lut_516_out;
    end
    endgenerate
    
    
    
    // LUT : 517
    wire [15:0] lut_517_table = 16'b1011111100000001;
    wire [3:0] lut_517_select = {
                             in_data[79],
                             in_data[231],
                             in_data[135],
                             in_data[21]};
    
    wire lut_517_out = lut_517_table[lut_517_select];
    
    generate
    if ( USE_REG ) begin : ff_517
        reg   lut_517_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_517_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_517_ff <= lut_517_out;
            end
        end
        
        assign out_data[517] = lut_517_ff;
    end
    else begin : no_ff_517
        assign out_data[517] = lut_517_out;
    end
    endgenerate
    
    
    
    // LUT : 518
    wire [15:0] lut_518_table = 16'b0010101010101010;
    wire [3:0] lut_518_select = {
                             in_data[146],
                             in_data[393],
                             in_data[34],
                             in_data[598]};
    
    wire lut_518_out = lut_518_table[lut_518_select];
    
    generate
    if ( USE_REG ) begin : ff_518
        reg   lut_518_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_518_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_518_ff <= lut_518_out;
            end
        end
        
        assign out_data[518] = lut_518_ff;
    end
    else begin : no_ff_518
        assign out_data[518] = lut_518_out;
    end
    endgenerate
    
    
    
    // LUT : 519
    wire [15:0] lut_519_table = 16'b0000001110111111;
    wire [3:0] lut_519_select = {
                             in_data[285],
                             in_data[19],
                             in_data[126],
                             in_data[526]};
    
    wire lut_519_out = lut_519_table[lut_519_select];
    
    generate
    if ( USE_REG ) begin : ff_519
        reg   lut_519_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_519_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_519_ff <= lut_519_out;
            end
        end
        
        assign out_data[519] = lut_519_ff;
    end
    else begin : no_ff_519
        assign out_data[519] = lut_519_out;
    end
    endgenerate
    
    
    
    // LUT : 520
    wire [15:0] lut_520_table = 16'b1011111110110000;
    wire [3:0] lut_520_select = {
                             in_data[560],
                             in_data[380],
                             in_data[354],
                             in_data[271]};
    
    wire lut_520_out = lut_520_table[lut_520_select];
    
    generate
    if ( USE_REG ) begin : ff_520
        reg   lut_520_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_520_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_520_ff <= lut_520_out;
            end
        end
        
        assign out_data[520] = lut_520_ff;
    end
    else begin : no_ff_520
        assign out_data[520] = lut_520_out;
    end
    endgenerate
    
    
    
    // LUT : 521
    wire [15:0] lut_521_table = 16'b1100111010001000;
    wire [3:0] lut_521_select = {
                             in_data[24],
                             in_data[430],
                             in_data[256],
                             in_data[501]};
    
    wire lut_521_out = lut_521_table[lut_521_select];
    
    generate
    if ( USE_REG ) begin : ff_521
        reg   lut_521_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_521_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_521_ff <= lut_521_out;
            end
        end
        
        assign out_data[521] = lut_521_ff;
    end
    else begin : no_ff_521
        assign out_data[521] = lut_521_out;
    end
    endgenerate
    
    
    
    // LUT : 522
    wire [15:0] lut_522_table = 16'b0000000011101111;
    wire [3:0] lut_522_select = {
                             in_data[429],
                             in_data[269],
                             in_data[571],
                             in_data[350]};
    
    wire lut_522_out = lut_522_table[lut_522_select];
    
    generate
    if ( USE_REG ) begin : ff_522
        reg   lut_522_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_522_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_522_ff <= lut_522_out;
            end
        end
        
        assign out_data[522] = lut_522_ff;
    end
    else begin : no_ff_522
        assign out_data[522] = lut_522_out;
    end
    endgenerate
    
    
    
    // LUT : 523
    wire [15:0] lut_523_table = 16'b0101000001010000;
    wire [3:0] lut_523_select = {
                             in_data[38],
                             in_data[523],
                             in_data[395],
                             in_data[463]};
    
    wire lut_523_out = lut_523_table[lut_523_select];
    
    generate
    if ( USE_REG ) begin : ff_523
        reg   lut_523_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_523_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_523_ff <= lut_523_out;
            end
        end
        
        assign out_data[523] = lut_523_ff;
    end
    else begin : no_ff_523
        assign out_data[523] = lut_523_out;
    end
    endgenerate
    
    
    
    // LUT : 524
    wire [15:0] lut_524_table = 16'b0000000001101111;
    wire [3:0] lut_524_select = {
                             in_data[440],
                             in_data[503],
                             in_data[74],
                             in_data[374]};
    
    wire lut_524_out = lut_524_table[lut_524_select];
    
    generate
    if ( USE_REG ) begin : ff_524
        reg   lut_524_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_524_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_524_ff <= lut_524_out;
            end
        end
        
        assign out_data[524] = lut_524_ff;
    end
    else begin : no_ff_524
        assign out_data[524] = lut_524_out;
    end
    endgenerate
    
    
    
    // LUT : 525
    wire [15:0] lut_525_table = 16'b0100010101011111;
    wire [3:0] lut_525_select = {
                             in_data[116],
                             in_data[376],
                             in_data[171],
                             in_data[635]};
    
    wire lut_525_out = lut_525_table[lut_525_select];
    
    generate
    if ( USE_REG ) begin : ff_525
        reg   lut_525_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_525_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_525_ff <= lut_525_out;
            end
        end
        
        assign out_data[525] = lut_525_ff;
    end
    else begin : no_ff_525
        assign out_data[525] = lut_525_out;
    end
    endgenerate
    
    
    
    // LUT : 526
    wire [15:0] lut_526_table = 16'b0100010001000100;
    wire [3:0] lut_526_select = {
                             in_data[92],
                             in_data[422],
                             in_data[114],
                             in_data[508]};
    
    wire lut_526_out = lut_526_table[lut_526_select];
    
    generate
    if ( USE_REG ) begin : ff_526
        reg   lut_526_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_526_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_526_ff <= lut_526_out;
            end
        end
        
        assign out_data[526] = lut_526_ff;
    end
    else begin : no_ff_526
        assign out_data[526] = lut_526_out;
    end
    endgenerate
    
    
    
    // LUT : 527
    wire [15:0] lut_527_table = 16'b1111111111011101;
    wire [3:0] lut_527_select = {
                             in_data[309],
                             in_data[3],
                             in_data[575],
                             in_data[442]};
    
    wire lut_527_out = lut_527_table[lut_527_select];
    
    generate
    if ( USE_REG ) begin : ff_527
        reg   lut_527_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_527_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_527_ff <= lut_527_out;
            end
        end
        
        assign out_data[527] = lut_527_ff;
    end
    else begin : no_ff_527
        assign out_data[527] = lut_527_out;
    end
    endgenerate
    
    
    
    // LUT : 528
    wire [15:0] lut_528_table = 16'b1010000010110010;
    wire [3:0] lut_528_select = {
                             in_data[110],
                             in_data[32],
                             in_data[154],
                             in_data[485]};
    
    wire lut_528_out = lut_528_table[lut_528_select];
    
    generate
    if ( USE_REG ) begin : ff_528
        reg   lut_528_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_528_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_528_ff <= lut_528_out;
            end
        end
        
        assign out_data[528] = lut_528_ff;
    end
    else begin : no_ff_528
        assign out_data[528] = lut_528_out;
    end
    endgenerate
    
    
    
    // LUT : 529
    wire [15:0] lut_529_table = 16'b1111111100000000;
    wire [3:0] lut_529_select = {
                             in_data[209],
                             in_data[330],
                             in_data[570],
                             in_data[213]};
    
    wire lut_529_out = lut_529_table[lut_529_select];
    
    generate
    if ( USE_REG ) begin : ff_529
        reg   lut_529_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_529_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_529_ff <= lut_529_out;
            end
        end
        
        assign out_data[529] = lut_529_ff;
    end
    else begin : no_ff_529
        assign out_data[529] = lut_529_out;
    end
    endgenerate
    
    
    
    // LUT : 530
    wire [15:0] lut_530_table = 16'b0010001010101010;
    wire [3:0] lut_530_select = {
                             in_data[315],
                             in_data[50],
                             in_data[275],
                             in_data[202]};
    
    wire lut_530_out = lut_530_table[lut_530_select];
    
    generate
    if ( USE_REG ) begin : ff_530
        reg   lut_530_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_530_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_530_ff <= lut_530_out;
            end
        end
        
        assign out_data[530] = lut_530_ff;
    end
    else begin : no_ff_530
        assign out_data[530] = lut_530_out;
    end
    endgenerate
    
    
    
    // LUT : 531
    wire [15:0] lut_531_table = 16'b1100000011101000;
    wire [3:0] lut_531_select = {
                             in_data[286],
                             in_data[122],
                             in_data[546],
                             in_data[351]};
    
    wire lut_531_out = lut_531_table[lut_531_select];
    
    generate
    if ( USE_REG ) begin : ff_531
        reg   lut_531_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_531_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_531_ff <= lut_531_out;
            end
        end
        
        assign out_data[531] = lut_531_ff;
    end
    else begin : no_ff_531
        assign out_data[531] = lut_531_out;
    end
    endgenerate
    
    
    
    // LUT : 532
    wire [15:0] lut_532_table = 16'b1101010011010101;
    wire [3:0] lut_532_select = {
                             in_data[131],
                             in_data[618],
                             in_data[208],
                             in_data[456]};
    
    wire lut_532_out = lut_532_table[lut_532_select];
    
    generate
    if ( USE_REG ) begin : ff_532
        reg   lut_532_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_532_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_532_ff <= lut_532_out;
            end
        end
        
        assign out_data[532] = lut_532_ff;
    end
    else begin : no_ff_532
        assign out_data[532] = lut_532_out;
    end
    endgenerate
    
    
    
    // LUT : 533
    wire [15:0] lut_533_table = 16'b0000000111001111;
    wire [3:0] lut_533_select = {
                             in_data[1],
                             in_data[466],
                             in_data[334],
                             in_data[359]};
    
    wire lut_533_out = lut_533_table[lut_533_select];
    
    generate
    if ( USE_REG ) begin : ff_533
        reg   lut_533_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_533_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_533_ff <= lut_533_out;
            end
        end
        
        assign out_data[533] = lut_533_ff;
    end
    else begin : no_ff_533
        assign out_data[533] = lut_533_out;
    end
    endgenerate
    
    
    
    // LUT : 534
    wire [15:0] lut_534_table = 16'b1010001010101010;
    wire [3:0] lut_534_select = {
                             in_data[207],
                             in_data[555],
                             in_data[600],
                             in_data[89]};
    
    wire lut_534_out = lut_534_table[lut_534_select];
    
    generate
    if ( USE_REG ) begin : ff_534
        reg   lut_534_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_534_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_534_ff <= lut_534_out;
            end
        end
        
        assign out_data[534] = lut_534_ff;
    end
    else begin : no_ff_534
        assign out_data[534] = lut_534_out;
    end
    endgenerate
    
    
    
    // LUT : 535
    wire [15:0] lut_535_table = 16'b0000100011101111;
    wire [3:0] lut_535_select = {
                             in_data[113],
                             in_data[587],
                             in_data[288],
                             in_data[121]};
    
    wire lut_535_out = lut_535_table[lut_535_select];
    
    generate
    if ( USE_REG ) begin : ff_535
        reg   lut_535_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_535_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_535_ff <= lut_535_out;
            end
        end
        
        assign out_data[535] = lut_535_ff;
    end
    else begin : no_ff_535
        assign out_data[535] = lut_535_out;
    end
    endgenerate
    
    
    
    // LUT : 536
    wire [15:0] lut_536_table = 16'b0000101100001011;
    wire [3:0] lut_536_select = {
                             in_data[270],
                             in_data[212],
                             in_data[347],
                             in_data[589]};
    
    wire lut_536_out = lut_536_table[lut_536_select];
    
    generate
    if ( USE_REG ) begin : ff_536
        reg   lut_536_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_536_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_536_ff <= lut_536_out;
            end
        end
        
        assign out_data[536] = lut_536_ff;
    end
    else begin : no_ff_536
        assign out_data[536] = lut_536_out;
    end
    endgenerate
    
    
    
    // LUT : 537
    wire [15:0] lut_537_table = 16'b0001111101001100;
    wire [3:0] lut_537_select = {
                             in_data[64],
                             in_data[424],
                             in_data[98],
                             in_data[167]};
    
    wire lut_537_out = lut_537_table[lut_537_select];
    
    generate
    if ( USE_REG ) begin : ff_537
        reg   lut_537_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_537_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_537_ff <= lut_537_out;
            end
        end
        
        assign out_data[537] = lut_537_ff;
    end
    else begin : no_ff_537
        assign out_data[537] = lut_537_out;
    end
    endgenerate
    
    
    
    // LUT : 538
    wire [15:0] lut_538_table = 16'b0001000011110000;
    wire [3:0] lut_538_select = {
                             in_data[336],
                             in_data[595],
                             in_data[406],
                             in_data[460]};
    
    wire lut_538_out = lut_538_table[lut_538_select];
    
    generate
    if ( USE_REG ) begin : ff_538
        reg   lut_538_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_538_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_538_ff <= lut_538_out;
            end
        end
        
        assign out_data[538] = lut_538_ff;
    end
    else begin : no_ff_538
        assign out_data[538] = lut_538_out;
    end
    endgenerate
    
    
    
    // LUT : 539
    wire [15:0] lut_539_table = 16'b0000010000001100;
    wire [3:0] lut_539_select = {
                             in_data[250],
                             in_data[631],
                             in_data[187],
                             in_data[450]};
    
    wire lut_539_out = lut_539_table[lut_539_select];
    
    generate
    if ( USE_REG ) begin : ff_539
        reg   lut_539_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_539_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_539_ff <= lut_539_out;
            end
        end
        
        assign out_data[539] = lut_539_ff;
    end
    else begin : no_ff_539
        assign out_data[539] = lut_539_out;
    end
    endgenerate
    
    
    
    // LUT : 540
    wire [15:0] lut_540_table = 16'b0101010011010100;
    wire [3:0] lut_540_select = {
                             in_data[47],
                             in_data[369],
                             in_data[509],
                             in_data[280]};
    
    wire lut_540_out = lut_540_table[lut_540_select];
    
    generate
    if ( USE_REG ) begin : ff_540
        reg   lut_540_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_540_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_540_ff <= lut_540_out;
            end
        end
        
        assign out_data[540] = lut_540_ff;
    end
    else begin : no_ff_540
        assign out_data[540] = lut_540_out;
    end
    endgenerate
    
    
    
    // LUT : 541
    wire [15:0] lut_541_table = 16'b1000100110000000;
    wire [3:0] lut_541_select = {
                             in_data[105],
                             in_data[473],
                             in_data[37],
                             in_data[175]};
    
    wire lut_541_out = lut_541_table[lut_541_select];
    
    generate
    if ( USE_REG ) begin : ff_541
        reg   lut_541_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_541_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_541_ff <= lut_541_out;
            end
        end
        
        assign out_data[541] = lut_541_ff;
    end
    else begin : no_ff_541
        assign out_data[541] = lut_541_out;
    end
    endgenerate
    
    
    
    // LUT : 542
    wire [15:0] lut_542_table = 16'b1111010111110101;
    wire [3:0] lut_542_select = {
                             in_data[408],
                             in_data[12],
                             in_data[353],
                             in_data[259]};
    
    wire lut_542_out = lut_542_table[lut_542_select];
    
    generate
    if ( USE_REG ) begin : ff_542
        reg   lut_542_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_542_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_542_ff <= lut_542_out;
            end
        end
        
        assign out_data[542] = lut_542_ff;
    end
    else begin : no_ff_542
        assign out_data[542] = lut_542_out;
    end
    endgenerate
    
    
    
    // LUT : 543
    wire [15:0] lut_543_table = 16'b1000000011001100;
    wire [3:0] lut_543_select = {
                             in_data[62],
                             in_data[470],
                             in_data[379],
                             in_data[124]};
    
    wire lut_543_out = lut_543_table[lut_543_select];
    
    generate
    if ( USE_REG ) begin : ff_543
        reg   lut_543_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_543_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_543_ff <= lut_543_out;
            end
        end
        
        assign out_data[543] = lut_543_ff;
    end
    else begin : no_ff_543
        assign out_data[543] = lut_543_out;
    end
    endgenerate
    
    
    
    // LUT : 544
    wire [15:0] lut_544_table = 16'b1111001101110101;
    wire [3:0] lut_544_select = {
                             in_data[561],
                             in_data[31],
                             in_data[317],
                             in_data[579]};
    
    wire lut_544_out = lut_544_table[lut_544_select];
    
    generate
    if ( USE_REG ) begin : ff_544
        reg   lut_544_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_544_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_544_ff <= lut_544_out;
            end
        end
        
        assign out_data[544] = lut_544_ff;
    end
    else begin : no_ff_544
        assign out_data[544] = lut_544_out;
    end
    endgenerate
    
    
    
    // LUT : 545
    wire [15:0] lut_545_table = 16'b0000111101001101;
    wire [3:0] lut_545_select = {
                             in_data[335],
                             in_data[273],
                             in_data[99],
                             in_data[211]};
    
    wire lut_545_out = lut_545_table[lut_545_select];
    
    generate
    if ( USE_REG ) begin : ff_545
        reg   lut_545_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_545_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_545_ff <= lut_545_out;
            end
        end
        
        assign out_data[545] = lut_545_ff;
    end
    else begin : no_ff_545
        assign out_data[545] = lut_545_out;
    end
    endgenerate
    
    
    
    // LUT : 546
    wire [15:0] lut_546_table = 16'b1111001000000010;
    wire [3:0] lut_546_select = {
                             in_data[582],
                             in_data[348],
                             in_data[100],
                             in_data[468]};
    
    wire lut_546_out = lut_546_table[lut_546_select];
    
    generate
    if ( USE_REG ) begin : ff_546
        reg   lut_546_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_546_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_546_ff <= lut_546_out;
            end
        end
        
        assign out_data[546] = lut_546_ff;
    end
    else begin : no_ff_546
        assign out_data[546] = lut_546_out;
    end
    endgenerate
    
    
    
    // LUT : 547
    wire [15:0] lut_547_table = 16'b1010111100001000;
    wire [3:0] lut_547_select = {
                             in_data[489],
                             in_data[569],
                             in_data[137],
                             in_data[198]};
    
    wire lut_547_out = lut_547_table[lut_547_select];
    
    generate
    if ( USE_REG ) begin : ff_547
        reg   lut_547_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_547_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_547_ff <= lut_547_out;
            end
        end
        
        assign out_data[547] = lut_547_ff;
    end
    else begin : no_ff_547
        assign out_data[547] = lut_547_out;
    end
    endgenerate
    
    
    
    // LUT : 548
    wire [15:0] lut_548_table = 16'b1111000011110001;
    wire [3:0] lut_548_select = {
                             in_data[253],
                             in_data[104],
                             in_data[342],
                             in_data[486]};
    
    wire lut_548_out = lut_548_table[lut_548_select];
    
    generate
    if ( USE_REG ) begin : ff_548
        reg   lut_548_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_548_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_548_ff <= lut_548_out;
            end
        end
        
        assign out_data[548] = lut_548_ff;
    end
    else begin : no_ff_548
        assign out_data[548] = lut_548_out;
    end
    endgenerate
    
    
    
    // LUT : 549
    wire [15:0] lut_549_table = 16'b1101010111111111;
    wire [3:0] lut_549_select = {
                             in_data[475],
                             in_data[293],
                             in_data[82],
                             in_data[610]};
    
    wire lut_549_out = lut_549_table[lut_549_select];
    
    generate
    if ( USE_REG ) begin : ff_549
        reg   lut_549_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_549_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_549_ff <= lut_549_out;
            end
        end
        
        assign out_data[549] = lut_549_ff;
    end
    else begin : no_ff_549
        assign out_data[549] = lut_549_out;
    end
    endgenerate
    
    
    
    // LUT : 550
    wire [15:0] lut_550_table = 16'b0001000001110000;
    wire [3:0] lut_550_select = {
                             in_data[195],
                             in_data[188],
                             in_data[563],
                             in_data[417]};
    
    wire lut_550_out = lut_550_table[lut_550_select];
    
    generate
    if ( USE_REG ) begin : ff_550
        reg   lut_550_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_550_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_550_ff <= lut_550_out;
            end
        end
        
        assign out_data[550] = lut_550_ff;
    end
    else begin : no_ff_550
        assign out_data[550] = lut_550_out;
    end
    endgenerate
    
    
    
    // LUT : 551
    wire [15:0] lut_551_table = 16'b0111111100000000;
    wire [3:0] lut_551_select = {
                             in_data[344],
                             in_data[479],
                             in_data[447],
                             in_data[320]};
    
    wire lut_551_out = lut_551_table[lut_551_select];
    
    generate
    if ( USE_REG ) begin : ff_551
        reg   lut_551_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_551_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_551_ff <= lut_551_out;
            end
        end
        
        assign out_data[551] = lut_551_ff;
    end
    else begin : no_ff_551
        assign out_data[551] = lut_551_out;
    end
    endgenerate
    
    
    
    // LUT : 552
    wire [15:0] lut_552_table = 16'b0000100010101011;
    wire [3:0] lut_552_select = {
                             in_data[243],
                             in_data[95],
                             in_data[318],
                             in_data[97]};
    
    wire lut_552_out = lut_552_table[lut_552_select];
    
    generate
    if ( USE_REG ) begin : ff_552
        reg   lut_552_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_552_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_552_ff <= lut_552_out;
            end
        end
        
        assign out_data[552] = lut_552_ff;
    end
    else begin : no_ff_552
        assign out_data[552] = lut_552_out;
    end
    endgenerate
    
    
    
    // LUT : 553
    wire [15:0] lut_553_table = 16'b0000101110101111;
    wire [3:0] lut_553_select = {
                             in_data[26],
                             in_data[13],
                             in_data[177],
                             in_data[107]};
    
    wire lut_553_out = lut_553_table[lut_553_select];
    
    generate
    if ( USE_REG ) begin : ff_553
        reg   lut_553_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_553_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_553_ff <= lut_553_out;
            end
        end
        
        assign out_data[553] = lut_553_ff;
    end
    else begin : no_ff_553
        assign out_data[553] = lut_553_out;
    end
    endgenerate
    
    
    
    // LUT : 554
    wire [15:0] lut_554_table = 16'b1010101011111111;
    wire [3:0] lut_554_select = {
                             in_data[36],
                             in_data[83],
                             in_data[229],
                             in_data[42]};
    
    wire lut_554_out = lut_554_table[lut_554_select];
    
    generate
    if ( USE_REG ) begin : ff_554
        reg   lut_554_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_554_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_554_ff <= lut_554_out;
            end
        end
        
        assign out_data[554] = lut_554_ff;
    end
    else begin : no_ff_554
        assign out_data[554] = lut_554_out;
    end
    endgenerate
    
    
    
    // LUT : 555
    wire [15:0] lut_555_table = 16'b0010000001010000;
    wire [3:0] lut_555_select = {
                             in_data[240],
                             in_data[559],
                             in_data[291],
                             in_data[597]};
    
    wire lut_555_out = lut_555_table[lut_555_select];
    
    generate
    if ( USE_REG ) begin : ff_555
        reg   lut_555_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_555_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_555_ff <= lut_555_out;
            end
        end
        
        assign out_data[555] = lut_555_ff;
    end
    else begin : no_ff_555
        assign out_data[555] = lut_555_out;
    end
    endgenerate
    
    
    
    // LUT : 556
    wire [15:0] lut_556_table = 16'b0011001011111010;
    wire [3:0] lut_556_select = {
                             in_data[40],
                             in_data[396],
                             in_data[609],
                             in_data[619]};
    
    wire lut_556_out = lut_556_table[lut_556_select];
    
    generate
    if ( USE_REG ) begin : ff_556
        reg   lut_556_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_556_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_556_ff <= lut_556_out;
            end
        end
        
        assign out_data[556] = lut_556_ff;
    end
    else begin : no_ff_556
        assign out_data[556] = lut_556_out;
    end
    endgenerate
    
    
    
    // LUT : 557
    wire [15:0] lut_557_table = 16'b0010001000111111;
    wire [3:0] lut_557_select = {
                             in_data[196],
                             in_data[605],
                             in_data[625],
                             in_data[482]};
    
    wire lut_557_out = lut_557_table[lut_557_select];
    
    generate
    if ( USE_REG ) begin : ff_557
        reg   lut_557_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_557_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_557_ff <= lut_557_out;
            end
        end
        
        assign out_data[557] = lut_557_ff;
    end
    else begin : no_ff_557
        assign out_data[557] = lut_557_out;
    end
    endgenerate
    
    
    
    // LUT : 558
    wire [15:0] lut_558_table = 16'b0011000011110011;
    wire [3:0] lut_558_select = {
                             in_data[515],
                             in_data[96],
                             in_data[169],
                             in_data[537]};
    
    wire lut_558_out = lut_558_table[lut_558_select];
    
    generate
    if ( USE_REG ) begin : ff_558
        reg   lut_558_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_558_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_558_ff <= lut_558_out;
            end
        end
        
        assign out_data[558] = lut_558_ff;
    end
    else begin : no_ff_558
        assign out_data[558] = lut_558_out;
    end
    endgenerate
    
    
    
    // LUT : 559
    wire [15:0] lut_559_table = 16'b1111011101110101;
    wire [3:0] lut_559_select = {
                             in_data[272],
                             in_data[7],
                             in_data[316],
                             in_data[592]};
    
    wire lut_559_out = lut_559_table[lut_559_select];
    
    generate
    if ( USE_REG ) begin : ff_559
        reg   lut_559_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_559_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_559_ff <= lut_559_out;
            end
        end
        
        assign out_data[559] = lut_559_ff;
    end
    else begin : no_ff_559
        assign out_data[559] = lut_559_out;
    end
    endgenerate
    
    
    
    // LUT : 560
    wire [15:0] lut_560_table = 16'b1100100011111111;
    wire [3:0] lut_560_select = {
                             in_data[329],
                             in_data[299],
                             in_data[49],
                             in_data[459]};
    
    wire lut_560_out = lut_560_table[lut_560_select];
    
    generate
    if ( USE_REG ) begin : ff_560
        reg   lut_560_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_560_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_560_ff <= lut_560_out;
            end
        end
        
        assign out_data[560] = lut_560_ff;
    end
    else begin : no_ff_560
        assign out_data[560] = lut_560_out;
    end
    endgenerate
    
    
    
    // LUT : 561
    wire [15:0] lut_561_table = 16'b1111111100100011;
    wire [3:0] lut_561_select = {
                             in_data[434],
                             in_data[54],
                             in_data[277],
                             in_data[517]};
    
    wire lut_561_out = lut_561_table[lut_561_select];
    
    generate
    if ( USE_REG ) begin : ff_561
        reg   lut_561_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_561_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_561_ff <= lut_561_out;
            end
        end
        
        assign out_data[561] = lut_561_ff;
    end
    else begin : no_ff_561
        assign out_data[561] = lut_561_out;
    end
    endgenerate
    
    
    
    // LUT : 562
    wire [15:0] lut_562_table = 16'b1011000011111010;
    wire [3:0] lut_562_select = {
                             in_data[580],
                             in_data[584],
                             in_data[65],
                             in_data[52]};
    
    wire lut_562_out = lut_562_table[lut_562_select];
    
    generate
    if ( USE_REG ) begin : ff_562
        reg   lut_562_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_562_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_562_ff <= lut_562_out;
            end
        end
        
        assign out_data[562] = lut_562_ff;
    end
    else begin : no_ff_562
        assign out_data[562] = lut_562_out;
    end
    endgenerate
    
    
    
    // LUT : 563
    wire [15:0] lut_563_table = 16'b0011001000110011;
    wire [3:0] lut_563_select = {
                             in_data[630],
                             in_data[585],
                             in_data[616],
                             in_data[77]};
    
    wire lut_563_out = lut_563_table[lut_563_select];
    
    generate
    if ( USE_REG ) begin : ff_563
        reg   lut_563_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_563_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_563_ff <= lut_563_out;
            end
        end
        
        assign out_data[563] = lut_563_ff;
    end
    else begin : no_ff_563
        assign out_data[563] = lut_563_out;
    end
    endgenerate
    
    
    
    // LUT : 564
    wire [15:0] lut_564_table = 16'b0001010100000001;
    wire [3:0] lut_564_select = {
                             in_data[67],
                             in_data[487],
                             in_data[18],
                             in_data[115]};
    
    wire lut_564_out = lut_564_table[lut_564_select];
    
    generate
    if ( USE_REG ) begin : ff_564
        reg   lut_564_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_564_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_564_ff <= lut_564_out;
            end
        end
        
        assign out_data[564] = lut_564_ff;
    end
    else begin : no_ff_564
        assign out_data[564] = lut_564_out;
    end
    endgenerate
    
    
    
    // LUT : 565
    wire [15:0] lut_565_table = 16'b0010001010111010;
    wire [3:0] lut_565_select = {
                             in_data[132],
                             in_data[70],
                             in_data[76],
                             in_data[588]};
    
    wire lut_565_out = lut_565_table[lut_565_select];
    
    generate
    if ( USE_REG ) begin : ff_565
        reg   lut_565_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_565_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_565_ff <= lut_565_out;
            end
        end
        
        assign out_data[565] = lut_565_ff;
    end
    else begin : no_ff_565
        assign out_data[565] = lut_565_out;
    end
    endgenerate
    
    
    
    // LUT : 566
    wire [15:0] lut_566_table = 16'b1101111011011111;
    wire [3:0] lut_566_select = {
                             in_data[224],
                             in_data[464],
                             in_data[282],
                             in_data[310]};
    
    wire lut_566_out = lut_566_table[lut_566_select];
    
    generate
    if ( USE_REG ) begin : ff_566
        reg   lut_566_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_566_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_566_ff <= lut_566_out;
            end
        end
        
        assign out_data[566] = lut_566_ff;
    end
    else begin : no_ff_566
        assign out_data[566] = lut_566_out;
    end
    endgenerate
    
    
    
    // LUT : 567
    wire [15:0] lut_567_table = 16'b0101111100001111;
    wire [3:0] lut_567_select = {
                             in_data[533],
                             in_data[136],
                             in_data[544],
                             in_data[254]};
    
    wire lut_567_out = lut_567_table[lut_567_select];
    
    generate
    if ( USE_REG ) begin : ff_567
        reg   lut_567_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_567_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_567_ff <= lut_567_out;
            end
        end
        
        assign out_data[567] = lut_567_ff;
    end
    else begin : no_ff_567
        assign out_data[567] = lut_567_out;
    end
    endgenerate
    
    
    
    // LUT : 568
    wire [15:0] lut_568_table = 16'b0100010011011111;
    wire [3:0] lut_568_select = {
                             in_data[409],
                             in_data[191],
                             in_data[203],
                             in_data[599]};
    
    wire lut_568_out = lut_568_table[lut_568_select];
    
    generate
    if ( USE_REG ) begin : ff_568
        reg   lut_568_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_568_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_568_ff <= lut_568_out;
            end
        end
        
        assign out_data[568] = lut_568_ff;
    end
    else begin : no_ff_568
        assign out_data[568] = lut_568_out;
    end
    endgenerate
    
    
    
    // LUT : 569
    wire [15:0] lut_569_table = 16'b1111110011111000;
    wire [3:0] lut_569_select = {
                             in_data[502],
                             in_data[433],
                             in_data[232],
                             in_data[25]};
    
    wire lut_569_out = lut_569_table[lut_569_select];
    
    generate
    if ( USE_REG ) begin : ff_569
        reg   lut_569_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_569_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_569_ff <= lut_569_out;
            end
        end
        
        assign out_data[569] = lut_569_ff;
    end
    else begin : no_ff_569
        assign out_data[569] = lut_569_out;
    end
    endgenerate
    
    
    
    // LUT : 570
    wire [15:0] lut_570_table = 16'b0011000010100000;
    wire [3:0] lut_570_select = {
                             in_data[357],
                             in_data[623],
                             in_data[390],
                             in_data[632]};
    
    wire lut_570_out = lut_570_table[lut_570_select];
    
    generate
    if ( USE_REG ) begin : ff_570
        reg   lut_570_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_570_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_570_ff <= lut_570_out;
            end
        end
        
        assign out_data[570] = lut_570_ff;
    end
    else begin : no_ff_570
        assign out_data[570] = lut_570_out;
    end
    endgenerate
    
    
    
    // LUT : 571
    wire [15:0] lut_571_table = 16'b0010000011111111;
    wire [3:0] lut_571_select = {
                             in_data[308],
                             in_data[452],
                             in_data[493],
                             in_data[483]};
    
    wire lut_571_out = lut_571_table[lut_571_select];
    
    generate
    if ( USE_REG ) begin : ff_571
        reg   lut_571_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_571_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_571_ff <= lut_571_out;
            end
        end
        
        assign out_data[571] = lut_571_ff;
    end
    else begin : no_ff_571
        assign out_data[571] = lut_571_out;
    end
    endgenerate
    
    
    
    // LUT : 572
    wire [15:0] lut_572_table = 16'b1111100011110000;
    wire [3:0] lut_572_select = {
                             in_data[614],
                             in_data[367],
                             in_data[119],
                             in_data[471]};
    
    wire lut_572_out = lut_572_table[lut_572_select];
    
    generate
    if ( USE_REG ) begin : ff_572
        reg   lut_572_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_572_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_572_ff <= lut_572_out;
            end
        end
        
        assign out_data[572] = lut_572_ff;
    end
    else begin : no_ff_572
        assign out_data[572] = lut_572_out;
    end
    endgenerate
    
    
    
    // LUT : 573
    wire [15:0] lut_573_table = 16'b0011000000110000;
    wire [3:0] lut_573_select = {
                             in_data[162],
                             in_data[613],
                             in_data[222],
                             in_data[248]};
    
    wire lut_573_out = lut_573_table[lut_573_select];
    
    generate
    if ( USE_REG ) begin : ff_573
        reg   lut_573_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_573_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_573_ff <= lut_573_out;
            end
        end
        
        assign out_data[573] = lut_573_ff;
    end
    else begin : no_ff_573
        assign out_data[573] = lut_573_out;
    end
    endgenerate
    
    
    
    // LUT : 574
    wire [15:0] lut_574_table = 16'b0010111100000000;
    wire [3:0] lut_574_select = {
                             in_data[276],
                             in_data[602],
                             in_data[166],
                             in_data[405]};
    
    wire lut_574_out = lut_574_table[lut_574_select];
    
    generate
    if ( USE_REG ) begin : ff_574
        reg   lut_574_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_574_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_574_ff <= lut_574_out;
            end
        end
        
        assign out_data[574] = lut_574_ff;
    end
    else begin : no_ff_574
        assign out_data[574] = lut_574_out;
    end
    endgenerate
    
    
    
    // LUT : 575
    wire [15:0] lut_575_table = 16'b0100010011111101;
    wire [3:0] lut_575_select = {
                             in_data[438],
                             in_data[45],
                             in_data[548],
                             in_data[492]};
    
    wire lut_575_out = lut_575_table[lut_575_select];
    
    generate
    if ( USE_REG ) begin : ff_575
        reg   lut_575_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_575_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_575_ff <= lut_575_out;
            end
        end
        
        assign out_data[575] = lut_575_ff;
    end
    else begin : no_ff_575
        assign out_data[575] = lut_575_out;
    end
    endgenerate
    
    
    
    // LUT : 576
    wire [15:0] lut_576_table = 16'b1101010111010101;
    wire [3:0] lut_576_select = {
                             in_data[633],
                             in_data[365],
                             in_data[193],
                             in_data[149]};
    
    wire lut_576_out = lut_576_table[lut_576_select];
    
    generate
    if ( USE_REG ) begin : ff_576
        reg   lut_576_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_576_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_576_ff <= lut_576_out;
            end
        end
        
        assign out_data[576] = lut_576_ff;
    end
    else begin : no_ff_576
        assign out_data[576] = lut_576_out;
    end
    endgenerate
    
    
    
    // LUT : 577
    wire [15:0] lut_577_table = 16'b1101110111011101;
    wire [3:0] lut_577_select = {
                             in_data[362],
                             in_data[120],
                             in_data[358],
                             in_data[205]};
    
    wire lut_577_out = lut_577_table[lut_577_select];
    
    generate
    if ( USE_REG ) begin : ff_577
        reg   lut_577_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_577_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_577_ff <= lut_577_out;
            end
        end
        
        assign out_data[577] = lut_577_ff;
    end
    else begin : no_ff_577
        assign out_data[577] = lut_577_out;
    end
    endgenerate
    
    
    
    // LUT : 578
    wire [15:0] lut_578_table = 16'b0101011101010111;
    wire [3:0] lut_578_select = {
                             in_data[9],
                             in_data[556],
                             in_data[201],
                             in_data[301]};
    
    wire lut_578_out = lut_578_table[lut_578_select];
    
    generate
    if ( USE_REG ) begin : ff_578
        reg   lut_578_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_578_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_578_ff <= lut_578_out;
            end
        end
        
        assign out_data[578] = lut_578_ff;
    end
    else begin : no_ff_578
        assign out_data[578] = lut_578_out;
    end
    endgenerate
    
    
    
    // LUT : 579
    wire [15:0] lut_579_table = 16'b0000000010111011;
    wire [3:0] lut_579_select = {
                             in_data[566],
                             in_data[455],
                             in_data[234],
                             in_data[152]};
    
    wire lut_579_out = lut_579_table[lut_579_select];
    
    generate
    if ( USE_REG ) begin : ff_579
        reg   lut_579_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_579_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_579_ff <= lut_579_out;
            end
        end
        
        assign out_data[579] = lut_579_ff;
    end
    else begin : no_ff_579
        assign out_data[579] = lut_579_out;
    end
    endgenerate
    
    
    
    // LUT : 580
    wire [15:0] lut_580_table = 16'b1111010001010000;
    wire [3:0] lut_580_select = {
                             in_data[314],
                             in_data[261],
                             in_data[22],
                             in_data[361]};
    
    wire lut_580_out = lut_580_table[lut_580_select];
    
    generate
    if ( USE_REG ) begin : ff_580
        reg   lut_580_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_580_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_580_ff <= lut_580_out;
            end
        end
        
        assign out_data[580] = lut_580_ff;
    end
    else begin : no_ff_580
        assign out_data[580] = lut_580_out;
    end
    endgenerate
    
    
    
    // LUT : 581
    wire [15:0] lut_581_table = 16'b0100110101011100;
    wire [3:0] lut_581_select = {
                             in_data[30],
                             in_data[27],
                             in_data[467],
                             in_data[128]};
    
    wire lut_581_out = lut_581_table[lut_581_select];
    
    generate
    if ( USE_REG ) begin : ff_581
        reg   lut_581_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_581_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_581_ff <= lut_581_out;
            end
        end
        
        assign out_data[581] = lut_581_ff;
    end
    else begin : no_ff_581
        assign out_data[581] = lut_581_out;
    end
    endgenerate
    
    
    
    // LUT : 582
    wire [15:0] lut_582_table = 16'b1101010101010100;
    wire [3:0] lut_582_select = {
                             in_data[245],
                             in_data[55],
                             in_data[304],
                             in_data[63]};
    
    wire lut_582_out = lut_582_table[lut_582_select];
    
    generate
    if ( USE_REG ) begin : ff_582
        reg   lut_582_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_582_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_582_ff <= lut_582_out;
            end
        end
        
        assign out_data[582] = lut_582_ff;
    end
    else begin : no_ff_582
        assign out_data[582] = lut_582_out;
    end
    endgenerate
    
    
    
    // LUT : 583
    wire [15:0] lut_583_table = 16'b1011111100101010;
    wire [3:0] lut_583_select = {
                             in_data[33],
                             in_data[477],
                             in_data[322],
                             in_data[525]};
    
    wire lut_583_out = lut_583_table[lut_583_select];
    
    generate
    if ( USE_REG ) begin : ff_583
        reg   lut_583_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_583_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_583_ff <= lut_583_out;
            end
        end
        
        assign out_data[583] = lut_583_ff;
    end
    else begin : no_ff_583
        assign out_data[583] = lut_583_out;
    end
    endgenerate
    
    
    
    // LUT : 584
    wire [15:0] lut_584_table = 16'b0000001100000011;
    wire [3:0] lut_584_select = {
                             in_data[303],
                             in_data[512],
                             in_data[217],
                             in_data[106]};
    
    wire lut_584_out = lut_584_table[lut_584_select];
    
    generate
    if ( USE_REG ) begin : ff_584
        reg   lut_584_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_584_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_584_ff <= lut_584_out;
            end
        end
        
        assign out_data[584] = lut_584_ff;
    end
    else begin : no_ff_584
        assign out_data[584] = lut_584_out;
    end
    endgenerate
    
    
    
    // LUT : 585
    wire [15:0] lut_585_table = 16'b1010101010101000;
    wire [3:0] lut_585_select = {
                             in_data[266],
                             in_data[494],
                             in_data[221],
                             in_data[530]};
    
    wire lut_585_out = lut_585_table[lut_585_select];
    
    generate
    if ( USE_REG ) begin : ff_585
        reg   lut_585_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_585_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_585_ff <= lut_585_out;
            end
        end
        
        assign out_data[585] = lut_585_ff;
    end
    else begin : no_ff_585
        assign out_data[585] = lut_585_out;
    end
    endgenerate
    
    
    
    // LUT : 586
    wire [15:0] lut_586_table = 16'b1100010011000100;
    wire [3:0] lut_586_select = {
                             in_data[325],
                             in_data[446],
                             in_data[506],
                             in_data[53]};
    
    wire lut_586_out = lut_586_table[lut_586_select];
    
    generate
    if ( USE_REG ) begin : ff_586
        reg   lut_586_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_586_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_586_ff <= lut_586_out;
            end
        end
        
        assign out_data[586] = lut_586_ff;
    end
    else begin : no_ff_586
        assign out_data[586] = lut_586_out;
    end
    endgenerate
    
    
    
    // LUT : 587
    wire [15:0] lut_587_table = 16'b1010001000100010;
    wire [3:0] lut_587_select = {
                             in_data[392],
                             in_data[23],
                             in_data[451],
                             in_data[58]};
    
    wire lut_587_out = lut_587_table[lut_587_select];
    
    generate
    if ( USE_REG ) begin : ff_587
        reg   lut_587_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_587_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_587_ff <= lut_587_out;
            end
        end
        
        assign out_data[587] = lut_587_ff;
    end
    else begin : no_ff_587
        assign out_data[587] = lut_587_out;
    end
    endgenerate
    
    
    
    // LUT : 588
    wire [15:0] lut_588_table = 16'b0111011100000101;
    wire [3:0] lut_588_select = {
                             in_data[535],
                             in_data[305],
                             in_data[192],
                             in_data[138]};
    
    wire lut_588_out = lut_588_table[lut_588_select];
    
    generate
    if ( USE_REG ) begin : ff_588
        reg   lut_588_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_588_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_588_ff <= lut_588_out;
            end
        end
        
        assign out_data[588] = lut_588_ff;
    end
    else begin : no_ff_588
        assign out_data[588] = lut_588_out;
    end
    endgenerate
    
    
    
    // LUT : 589
    wire [15:0] lut_589_table = 16'b0010001000110011;
    wire [3:0] lut_589_select = {
                             in_data[182],
                             in_data[608],
                             in_data[534],
                             in_data[427]};
    
    wire lut_589_out = lut_589_table[lut_589_select];
    
    generate
    if ( USE_REG ) begin : ff_589
        reg   lut_589_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_589_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_589_ff <= lut_589_out;
            end
        end
        
        assign out_data[589] = lut_589_ff;
    end
    else begin : no_ff_589
        assign out_data[589] = lut_589_out;
    end
    endgenerate
    
    
    
    // LUT : 590
    wire [15:0] lut_590_table = 16'b0000010001010101;
    wire [3:0] lut_590_select = {
                             in_data[225],
                             in_data[284],
                             in_data[394],
                             in_data[524]};
    
    wire lut_590_out = lut_590_table[lut_590_select];
    
    generate
    if ( USE_REG ) begin : ff_590
        reg   lut_590_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_590_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_590_ff <= lut_590_out;
            end
        end
        
        assign out_data[590] = lut_590_ff;
    end
    else begin : no_ff_590
        assign out_data[590] = lut_590_out;
    end
    endgenerate
    
    
    
    // LUT : 591
    wire [15:0] lut_591_table = 16'b0001000100010111;
    wire [3:0] lut_591_select = {
                             in_data[326],
                             in_data[345],
                             in_data[421],
                             in_data[289]};
    
    wire lut_591_out = lut_591_table[lut_591_select];
    
    generate
    if ( USE_REG ) begin : ff_591
        reg   lut_591_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_591_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_591_ff <= lut_591_out;
            end
        end
        
        assign out_data[591] = lut_591_ff;
    end
    else begin : no_ff_591
        assign out_data[591] = lut_591_out;
    end
    endgenerate
    
    
    
    // LUT : 592
    wire [15:0] lut_592_table = 16'b0000000000010111;
    wire [3:0] lut_592_select = {
                             in_data[536],
                             in_data[144],
                             in_data[60],
                             in_data[622]};
    
    wire lut_592_out = lut_592_table[lut_592_select];
    
    generate
    if ( USE_REG ) begin : ff_592
        reg   lut_592_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_592_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_592_ff <= lut_592_out;
            end
        end
        
        assign out_data[592] = lut_592_ff;
    end
    else begin : no_ff_592
        assign out_data[592] = lut_592_out;
    end
    endgenerate
    
    
    
    // LUT : 593
    wire [15:0] lut_593_table = 16'b0000011100010101;
    wire [3:0] lut_593_select = {
                             in_data[539],
                             in_data[183],
                             in_data[435],
                             in_data[577]};
    
    wire lut_593_out = lut_593_table[lut_593_select];
    
    generate
    if ( USE_REG ) begin : ff_593
        reg   lut_593_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_593_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_593_ff <= lut_593_out;
            end
        end
        
        assign out_data[593] = lut_593_ff;
    end
    else begin : no_ff_593
        assign out_data[593] = lut_593_out;
    end
    endgenerate
    
    
    
    // LUT : 594
    wire [15:0] lut_594_table = 16'b0001000001010101;
    wire [3:0] lut_594_select = {
                             in_data[84],
                             in_data[403],
                             in_data[313],
                             in_data[385]};
    
    wire lut_594_out = lut_594_table[lut_594_select];
    
    generate
    if ( USE_REG ) begin : ff_594
        reg   lut_594_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_594_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_594_ff <= lut_594_out;
            end
        end
        
        assign out_data[594] = lut_594_ff;
    end
    else begin : no_ff_594
        assign out_data[594] = lut_594_out;
    end
    endgenerate
    
    
    
    // LUT : 595
    wire [15:0] lut_595_table = 16'b0010000010110010;
    wire [3:0] lut_595_select = {
                             in_data[527],
                             in_data[415],
                             in_data[543],
                             in_data[499]};
    
    wire lut_595_out = lut_595_table[lut_595_select];
    
    generate
    if ( USE_REG ) begin : ff_595
        reg   lut_595_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_595_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_595_ff <= lut_595_out;
            end
        end
        
        assign out_data[595] = lut_595_ff;
    end
    else begin : no_ff_595
        assign out_data[595] = lut_595_out;
    end
    endgenerate
    
    
    
    // LUT : 596
    wire [15:0] lut_596_table = 16'b1000110010001110;
    wire [3:0] lut_596_select = {
                             in_data[397],
                             in_data[75],
                             in_data[287],
                             in_data[71]};
    
    wire lut_596_out = lut_596_table[lut_596_select];
    
    generate
    if ( USE_REG ) begin : ff_596
        reg   lut_596_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_596_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_596_ff <= lut_596_out;
            end
        end
        
        assign out_data[596] = lut_596_ff;
    end
    else begin : no_ff_596
        assign out_data[596] = lut_596_out;
    end
    endgenerate
    
    
    
    // LUT : 597
    wire [15:0] lut_597_table = 16'b0000000001001111;
    wire [3:0] lut_597_select = {
                             in_data[510],
                             in_data[457],
                             in_data[189],
                             in_data[168]};
    
    wire lut_597_out = lut_597_table[lut_597_select];
    
    generate
    if ( USE_REG ) begin : ff_597
        reg   lut_597_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_597_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_597_ff <= lut_597_out;
            end
        end
        
        assign out_data[597] = lut_597_ff;
    end
    else begin : no_ff_597
        assign out_data[597] = lut_597_out;
    end
    endgenerate
    
    
    
    // LUT : 598
    wire [15:0] lut_598_table = 16'b0101000011010101;
    wire [3:0] lut_598_select = {
                             in_data[158],
                             in_data[352],
                             in_data[449],
                             in_data[164]};
    
    wire lut_598_out = lut_598_table[lut_598_select];
    
    generate
    if ( USE_REG ) begin : ff_598
        reg   lut_598_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_598_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_598_ff <= lut_598_out;
            end
        end
        
        assign out_data[598] = lut_598_ff;
    end
    else begin : no_ff_598
        assign out_data[598] = lut_598_out;
    end
    endgenerate
    
    
    
    // LUT : 599
    wire [15:0] lut_599_table = 16'b0001010100010001;
    wire [3:0] lut_599_select = {
                             in_data[431],
                             in_data[165],
                             in_data[549],
                             in_data[176]};
    
    wire lut_599_out = lut_599_table[lut_599_select];
    
    generate
    if ( USE_REG ) begin : ff_599
        reg   lut_599_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_599_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_599_ff <= lut_599_out;
            end
        end
        
        assign out_data[599] = lut_599_ff;
    end
    else begin : no_ff_599
        assign out_data[599] = lut_599_out;
    end
    endgenerate
    
    
    
    // LUT : 600
    wire [15:0] lut_600_table = 16'b1100111111111010;
    wire [3:0] lut_600_select = {
                             in_data[279],
                             in_data[495],
                             in_data[377],
                             in_data[491]};
    
    wire lut_600_out = lut_600_table[lut_600_select];
    
    generate
    if ( USE_REG ) begin : ff_600
        reg   lut_600_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_600_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_600_ff <= lut_600_out;
            end
        end
        
        assign out_data[600] = lut_600_ff;
    end
    else begin : no_ff_600
        assign out_data[600] = lut_600_out;
    end
    endgenerate
    
    
    
    // LUT : 601
    wire [15:0] lut_601_table = 16'b1110110011101000;
    wire [3:0] lut_601_select = {
                             in_data[8],
                             in_data[87],
                             in_data[480],
                             in_data[338]};
    
    wire lut_601_out = lut_601_table[lut_601_select];
    
    generate
    if ( USE_REG ) begin : ff_601
        reg   lut_601_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_601_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_601_ff <= lut_601_out;
            end
        end
        
        assign out_data[601] = lut_601_ff;
    end
    else begin : no_ff_601
        assign out_data[601] = lut_601_out;
    end
    endgenerate
    
    
    
    // LUT : 602
    wire [15:0] lut_602_table = 16'b1111000011111100;
    wire [3:0] lut_602_select = {
                             in_data[505],
                             in_data[565],
                             in_data[391],
                             in_data[43]};
    
    wire lut_602_out = lut_602_table[lut_602_select];
    
    generate
    if ( USE_REG ) begin : ff_602
        reg   lut_602_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_602_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_602_ff <= lut_602_out;
            end
        end
        
        assign out_data[602] = lut_602_ff;
    end
    else begin : no_ff_602
        assign out_data[602] = lut_602_out;
    end
    endgenerate
    
    
    
    // LUT : 603
    wire [15:0] lut_603_table = 16'b1111001010110010;
    wire [3:0] lut_603_select = {
                             in_data[545],
                             in_data[156],
                             in_data[159],
                             in_data[603]};
    
    wire lut_603_out = lut_603_table[lut_603_select];
    
    generate
    if ( USE_REG ) begin : ff_603
        reg   lut_603_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_603_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_603_ff <= lut_603_out;
            end
        end
        
        assign out_data[603] = lut_603_ff;
    end
    else begin : no_ff_603
        assign out_data[603] = lut_603_out;
    end
    endgenerate
    
    
    
    // LUT : 604
    wire [15:0] lut_604_table = 16'b1100111100001100;
    wire [3:0] lut_604_select = {
                             in_data[214],
                             in_data[20],
                             in_data[139],
                             in_data[219]};
    
    wire lut_604_out = lut_604_table[lut_604_select];
    
    generate
    if ( USE_REG ) begin : ff_604
        reg   lut_604_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_604_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_604_ff <= lut_604_out;
            end
        end
        
        assign out_data[604] = lut_604_ff;
    end
    else begin : no_ff_604
        assign out_data[604] = lut_604_out;
    end
    endgenerate
    
    
    
    // LUT : 605
    wire [15:0] lut_605_table = 16'b1111110111110101;
    wire [3:0] lut_605_select = {
                             in_data[111],
                             in_data[161],
                             in_data[606],
                             in_data[11]};
    
    wire lut_605_out = lut_605_table[lut_605_select];
    
    generate
    if ( USE_REG ) begin : ff_605
        reg   lut_605_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_605_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_605_ff <= lut_605_out;
            end
        end
        
        assign out_data[605] = lut_605_ff;
    end
    else begin : no_ff_605
        assign out_data[605] = lut_605_out;
    end
    endgenerate
    
    
    
    // LUT : 606
    wire [15:0] lut_606_table = 16'b1111101010000000;
    wire [3:0] lut_606_select = {
                             in_data[102],
                             in_data[295],
                             in_data[568],
                             in_data[615]};
    
    wire lut_606_out = lut_606_table[lut_606_select];
    
    generate
    if ( USE_REG ) begin : ff_606
        reg   lut_606_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_606_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_606_ff <= lut_606_out;
            end
        end
        
        assign out_data[606] = lut_606_ff;
    end
    else begin : no_ff_606
        assign out_data[606] = lut_606_out;
    end
    endgenerate
    
    
    
    // LUT : 607
    wire [15:0] lut_607_table = 16'b1111001100100000;
    wire [3:0] lut_607_select = {
                             in_data[147],
                             in_data[381],
                             in_data[339],
                             in_data[436]};
    
    wire lut_607_out = lut_607_table[lut_607_select];
    
    generate
    if ( USE_REG ) begin : ff_607
        reg   lut_607_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_607_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_607_ff <= lut_607_out;
            end
        end
        
        assign out_data[607] = lut_607_ff;
    end
    else begin : no_ff_607
        assign out_data[607] = lut_607_out;
    end
    endgenerate
    
    
    
    // LUT : 608
    wire [15:0] lut_608_table = 16'b1010000011101110;
    wire [3:0] lut_608_select = {
                             in_data[230],
                             in_data[260],
                             in_data[108],
                             in_data[94]};
    
    wire lut_608_out = lut_608_table[lut_608_select];
    
    generate
    if ( USE_REG ) begin : ff_608
        reg   lut_608_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_608_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_608_ff <= lut_608_out;
            end
        end
        
        assign out_data[608] = lut_608_ff;
    end
    else begin : no_ff_608
        assign out_data[608] = lut_608_out;
    end
    endgenerate
    
    
    
    // LUT : 609
    wire [15:0] lut_609_table = 16'b1101000011110100;
    wire [3:0] lut_609_select = {
                             in_data[611],
                             in_data[233],
                             in_data[593],
                             in_data[364]};
    
    wire lut_609_out = lut_609_table[lut_609_select];
    
    generate
    if ( USE_REG ) begin : ff_609
        reg   lut_609_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_609_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_609_ff <= lut_609_out;
            end
        end
        
        assign out_data[609] = lut_609_ff;
    end
    else begin : no_ff_609
        assign out_data[609] = lut_609_out;
    end
    endgenerate
    
    
    
    // LUT : 610
    wire [15:0] lut_610_table = 16'b0000001011111011;
    wire [3:0] lut_610_select = {
                             in_data[578],
                             in_data[197],
                             in_data[312],
                             in_data[514]};
    
    wire lut_610_out = lut_610_table[lut_610_select];
    
    generate
    if ( USE_REG ) begin : ff_610
        reg   lut_610_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_610_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_610_ff <= lut_610_out;
            end
        end
        
        assign out_data[610] = lut_610_ff;
    end
    else begin : no_ff_610
        assign out_data[610] = lut_610_out;
    end
    endgenerate
    
    
    
    // LUT : 611
    wire [15:0] lut_611_table = 16'b0010001110110011;
    wire [3:0] lut_611_select = {
                             in_data[319],
                             in_data[226],
                             in_data[636],
                             in_data[244]};
    
    wire lut_611_out = lut_611_table[lut_611_select];
    
    generate
    if ( USE_REG ) begin : ff_611
        reg   lut_611_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_611_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_611_ff <= lut_611_out;
            end
        end
        
        assign out_data[611] = lut_611_ff;
    end
    else begin : no_ff_611
        assign out_data[611] = lut_611_out;
    end
    endgenerate
    
    
    
    // LUT : 612
    wire [15:0] lut_612_table = 16'b1000110110001100;
    wire [3:0] lut_612_select = {
                             in_data[574],
                             in_data[29],
                             in_data[306],
                             in_data[551]};
    
    wire lut_612_out = lut_612_table[lut_612_select];
    
    generate
    if ( USE_REG ) begin : ff_612
        reg   lut_612_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_612_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_612_ff <= lut_612_out;
            end
        end
        
        assign out_data[612] = lut_612_ff;
    end
    else begin : no_ff_612
        assign out_data[612] = lut_612_out;
    end
    endgenerate
    
    
    
    // LUT : 613
    wire [15:0] lut_613_table = 16'b1010100011101010;
    wire [3:0] lut_613_select = {
                             in_data[437],
                             in_data[404],
                             in_data[343],
                             in_data[86]};
    
    wire lut_613_out = lut_613_table[lut_613_select];
    
    generate
    if ( USE_REG ) begin : ff_613
        reg   lut_613_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_613_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_613_ff <= lut_613_out;
            end
        end
        
        assign out_data[613] = lut_613_ff;
    end
    else begin : no_ff_613
        assign out_data[613] = lut_613_out;
    end
    endgenerate
    
    
    
    // LUT : 614
    wire [15:0] lut_614_table = 16'b1100110000000000;
    wire [3:0] lut_614_select = {
                             in_data[454],
                             in_data[194],
                             in_data[160],
                             in_data[507]};
    
    wire lut_614_out = lut_614_table[lut_614_select];
    
    generate
    if ( USE_REG ) begin : ff_614
        reg   lut_614_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_614_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_614_ff <= lut_614_out;
            end
        end
        
        assign out_data[614] = lut_614_ff;
    end
    else begin : no_ff_614
        assign out_data[614] = lut_614_out;
    end
    endgenerate
    
    
    
    // LUT : 615
    wire [15:0] lut_615_table = 16'b1000111010111111;
    wire [3:0] lut_615_select = {
                             in_data[553],
                             in_data[81],
                             in_data[93],
                             in_data[423]};
    
    wire lut_615_out = lut_615_table[lut_615_select];
    
    generate
    if ( USE_REG ) begin : ff_615
        reg   lut_615_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_615_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_615_ff <= lut_615_out;
            end
        end
        
        assign out_data[615] = lut_615_ff;
    end
    else begin : no_ff_615
        assign out_data[615] = lut_615_out;
    end
    endgenerate
    
    
    
    // LUT : 616
    wire [15:0] lut_616_table = 16'b1011100111110100;
    wire [3:0] lut_616_select = {
                             in_data[418],
                             in_data[383],
                             in_data[583],
                             in_data[141]};
    
    wire lut_616_out = lut_616_table[lut_616_select];
    
    generate
    if ( USE_REG ) begin : ff_616
        reg   lut_616_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_616_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_616_ff <= lut_616_out;
            end
        end
        
        assign out_data[616] = lut_616_ff;
    end
    else begin : no_ff_616
        assign out_data[616] = lut_616_out;
    end
    endgenerate
    
    
    
    // LUT : 617
    wire [15:0] lut_617_table = 16'b1101110101010100;
    wire [3:0] lut_617_select = {
                             in_data[298],
                             in_data[15],
                             in_data[621],
                             in_data[220]};
    
    wire lut_617_out = lut_617_table[lut_617_select];
    
    generate
    if ( USE_REG ) begin : ff_617
        reg   lut_617_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_617_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_617_ff <= lut_617_out;
            end
        end
        
        assign out_data[617] = lut_617_ff;
    end
    else begin : no_ff_617
        assign out_data[617] = lut_617_out;
    end
    endgenerate
    
    
    
    // LUT : 618
    wire [15:0] lut_618_table = 16'b1010101110100011;
    wire [3:0] lut_618_select = {
                             in_data[637],
                             in_data[66],
                             in_data[432],
                             in_data[627]};
    
    wire lut_618_out = lut_618_table[lut_618_select];
    
    generate
    if ( USE_REG ) begin : ff_618
        reg   lut_618_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_618_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_618_ff <= lut_618_out;
            end
        end
        
        assign out_data[618] = lut_618_ff;
    end
    else begin : no_ff_618
        assign out_data[618] = lut_618_out;
    end
    endgenerate
    
    
    
    // LUT : 619
    wire [15:0] lut_619_table = 16'b1111001100000000;
    wire [3:0] lut_619_select = {
                             in_data[179],
                             in_data[206],
                             in_data[371],
                             in_data[163]};
    
    wire lut_619_out = lut_619_table[lut_619_select];
    
    generate
    if ( USE_REG ) begin : ff_619
        reg   lut_619_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_619_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_619_ff <= lut_619_out;
            end
        end
        
        assign out_data[619] = lut_619_ff;
    end
    else begin : no_ff_619
        assign out_data[619] = lut_619_out;
    end
    endgenerate
    
    
    
    // LUT : 620
    wire [15:0] lut_620_table = 16'b1110100011111110;
    wire [3:0] lut_620_select = {
                             in_data[378],
                             in_data[529],
                             in_data[400],
                             in_data[497]};
    
    wire lut_620_out = lut_620_table[lut_620_select];
    
    generate
    if ( USE_REG ) begin : ff_620
        reg   lut_620_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_620_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_620_ff <= lut_620_out;
            end
        end
        
        assign out_data[620] = lut_620_ff;
    end
    else begin : no_ff_620
        assign out_data[620] = lut_620_out;
    end
    endgenerate
    
    
    
    // LUT : 621
    wire [15:0] lut_621_table = 16'b0011011101110011;
    wire [3:0] lut_621_select = {
                             in_data[458],
                             in_data[384],
                             in_data[370],
                             in_data[184]};
    
    wire lut_621_out = lut_621_table[lut_621_select];
    
    generate
    if ( USE_REG ) begin : ff_621
        reg   lut_621_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_621_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_621_ff <= lut_621_out;
            end
        end
        
        assign out_data[621] = lut_621_ff;
    end
    else begin : no_ff_621
        assign out_data[621] = lut_621_out;
    end
    endgenerate
    
    
    
    // LUT : 622
    wire [15:0] lut_622_table = 16'b0000010000101111;
    wire [3:0] lut_622_select = {
                             in_data[210],
                             in_data[56],
                             in_data[69],
                             in_data[518]};
    
    wire lut_622_out = lut_622_table[lut_622_select];
    
    generate
    if ( USE_REG ) begin : ff_622
        reg   lut_622_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_622_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_622_ff <= lut_622_out;
            end
        end
        
        assign out_data[622] = lut_622_ff;
    end
    else begin : no_ff_622
        assign out_data[622] = lut_622_out;
    end
    endgenerate
    
    
    
    // LUT : 623
    wire [15:0] lut_623_table = 16'b1101110101010100;
    wire [3:0] lut_623_select = {
                             in_data[469],
                             in_data[150],
                             in_data[117],
                             in_data[247]};
    
    wire lut_623_out = lut_623_table[lut_623_select];
    
    generate
    if ( USE_REG ) begin : ff_623
        reg   lut_623_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_623_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_623_ff <= lut_623_out;
            end
        end
        
        assign out_data[623] = lut_623_ff;
    end
    else begin : no_ff_623
        assign out_data[623] = lut_623_out;
    end
    endgenerate
    
    
    
    // LUT : 624
    wire [15:0] lut_624_table = 16'b1010101110111011;
    wire [3:0] lut_624_select = {
                             in_data[538],
                             in_data[181],
                             in_data[16],
                             in_data[281]};
    
    wire lut_624_out = lut_624_table[lut_624_select];
    
    generate
    if ( USE_REG ) begin : ff_624
        reg   lut_624_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_624_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_624_ff <= lut_624_out;
            end
        end
        
        assign out_data[624] = lut_624_ff;
    end
    else begin : no_ff_624
        assign out_data[624] = lut_624_out;
    end
    endgenerate
    
    
    
    // LUT : 625
    wire [15:0] lut_625_table = 16'b0101010100000000;
    wire [3:0] lut_625_select = {
                             in_data[257],
                             in_data[242],
                             in_data[237],
                             in_data[216]};
    
    wire lut_625_out = lut_625_table[lut_625_select];
    
    generate
    if ( USE_REG ) begin : ff_625
        reg   lut_625_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_625_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_625_ff <= lut_625_out;
            end
        end
        
        assign out_data[625] = lut_625_ff;
    end
    else begin : no_ff_625
        assign out_data[625] = lut_625_out;
    end
    endgenerate
    
    
    
    // LUT : 626
    wire [15:0] lut_626_table = 16'b0011011100000000;
    wire [3:0] lut_626_select = {
                             in_data[265],
                             in_data[341],
                             in_data[17],
                             in_data[366]};
    
    wire lut_626_out = lut_626_table[lut_626_select];
    
    generate
    if ( USE_REG ) begin : ff_626
        reg   lut_626_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_626_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_626_ff <= lut_626_out;
            end
        end
        
        assign out_data[626] = lut_626_ff;
    end
    else begin : no_ff_626
        assign out_data[626] = lut_626_out;
    end
    endgenerate
    
    
    
    // LUT : 627
    wire [15:0] lut_627_table = 16'b0000000001001101;
    wire [3:0] lut_627_select = {
                             in_data[476],
                             in_data[241],
                             in_data[48],
                             in_data[331]};
    
    wire lut_627_out = lut_627_table[lut_627_select];
    
    generate
    if ( USE_REG ) begin : ff_627
        reg   lut_627_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_627_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_627_ff <= lut_627_out;
            end
        end
        
        assign out_data[627] = lut_627_ff;
    end
    else begin : no_ff_627
        assign out_data[627] = lut_627_out;
    end
    endgenerate
    
    
    
    // LUT : 628
    wire [15:0] lut_628_table = 16'b0100010001010100;
    wire [3:0] lut_628_select = {
                             in_data[51],
                             in_data[356],
                             in_data[57],
                             in_data[324]};
    
    wire lut_628_out = lut_628_table[lut_628_select];
    
    generate
    if ( USE_REG ) begin : ff_628
        reg   lut_628_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_628_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_628_ff <= lut_628_out;
            end
        end
        
        assign out_data[628] = lut_628_ff;
    end
    else begin : no_ff_628
        assign out_data[628] = lut_628_out;
    end
    endgenerate
    
    
    
    // LUT : 629
    wire [15:0] lut_629_table = 16'b1111111100000000;
    wire [3:0] lut_629_select = {
                             in_data[401],
                             in_data[528],
                             in_data[620],
                             in_data[412]};
    
    wire lut_629_out = lut_629_table[lut_629_select];
    
    generate
    if ( USE_REG ) begin : ff_629
        reg   lut_629_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_629_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_629_ff <= lut_629_out;
            end
        end
        
        assign out_data[629] = lut_629_ff;
    end
    else begin : no_ff_629
        assign out_data[629] = lut_629_out;
    end
    endgenerate
    
    
    
    // LUT : 630
    wire [15:0] lut_630_table = 16'b1100111100001000;
    wire [3:0] lut_630_select = {
                             in_data[488],
                             in_data[4],
                             in_data[541],
                             in_data[590]};
    
    wire lut_630_out = lut_630_table[lut_630_select];
    
    generate
    if ( USE_REG ) begin : ff_630
        reg   lut_630_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_630_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_630_ff <= lut_630_out;
            end
        end
        
        assign out_data[630] = lut_630_ff;
    end
    else begin : no_ff_630
        assign out_data[630] = lut_630_out;
    end
    endgenerate
    
    
    
    // LUT : 631
    wire [15:0] lut_631_table = 16'b0000001000011111;
    wire [3:0] lut_631_select = {
                             in_data[581],
                             in_data[80],
                             in_data[388],
                             in_data[386]};
    
    wire lut_631_out = lut_631_table[lut_631_select];
    
    generate
    if ( USE_REG ) begin : ff_631
        reg   lut_631_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_631_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_631_ff <= lut_631_out;
            end
        end
        
        assign out_data[631] = lut_631_ff;
    end
    else begin : no_ff_631
        assign out_data[631] = lut_631_out;
    end
    endgenerate
    
    
    
    // LUT : 632
    wire [15:0] lut_632_table = 16'b0000110011001111;
    wire [3:0] lut_632_select = {
                             in_data[123],
                             in_data[173],
                             in_data[594],
                             in_data[490]};
    
    wire lut_632_out = lut_632_table[lut_632_select];
    
    generate
    if ( USE_REG ) begin : ff_632
        reg   lut_632_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_632_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_632_ff <= lut_632_out;
            end
        end
        
        assign out_data[632] = lut_632_ff;
    end
    else begin : no_ff_632
        assign out_data[632] = lut_632_out;
    end
    endgenerate
    
    
    
    // LUT : 633
    wire [15:0] lut_633_table = 16'b1110111011101110;
    wire [3:0] lut_633_select = {
                             in_data[252],
                             in_data[498],
                             in_data[307],
                             in_data[215]};
    
    wire lut_633_out = lut_633_table[lut_633_select];
    
    generate
    if ( USE_REG ) begin : ff_633
        reg   lut_633_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_633_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_633_ff <= lut_633_out;
            end
        end
        
        assign out_data[633] = lut_633_ff;
    end
    else begin : no_ff_633
        assign out_data[633] = lut_633_out;
    end
    endgenerate
    
    
    
    // LUT : 634
    wire [15:0] lut_634_table = 16'b1111101110110000;
    wire [3:0] lut_634_select = {
                             in_data[607],
                             in_data[186],
                             in_data[327],
                             in_data[372]};
    
    wire lut_634_out = lut_634_table[lut_634_select];
    
    generate
    if ( USE_REG ) begin : ff_634
        reg   lut_634_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_634_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_634_ff <= lut_634_out;
            end
        end
        
        assign out_data[634] = lut_634_ff;
    end
    else begin : no_ff_634
        assign out_data[634] = lut_634_out;
    end
    endgenerate
    
    
    
    // LUT : 635
    wire [15:0] lut_635_table = 16'b1010001010101010;
    wire [3:0] lut_635_select = {
                             in_data[398],
                             in_data[311],
                             in_data[612],
                             in_data[441]};
    
    wire lut_635_out = lut_635_table[lut_635_select];
    
    generate
    if ( USE_REG ) begin : ff_635
        reg   lut_635_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_635_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_635_ff <= lut_635_out;
            end
        end
        
        assign out_data[635] = lut_635_ff;
    end
    else begin : no_ff_635
        assign out_data[635] = lut_635_out;
    end
    endgenerate
    
    
    
    // LUT : 636
    wire [15:0] lut_636_table = 16'b1010001011101010;
    wire [3:0] lut_636_select = {
                             in_data[278],
                             in_data[85],
                             in_data[382],
                             in_data[474]};
    
    wire lut_636_out = lut_636_table[lut_636_select];
    
    generate
    if ( USE_REG ) begin : ff_636
        reg   lut_636_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_636_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_636_ff <= lut_636_out;
            end
        end
        
        assign out_data[636] = lut_636_ff;
    end
    else begin : no_ff_636
        assign out_data[636] = lut_636_out;
    end
    endgenerate
    
    
    
    // LUT : 637
    wire [15:0] lut_637_table = 16'b0010111111101110;
    wire [3:0] lut_637_select = {
                             in_data[263],
                             in_data[500],
                             in_data[218],
                             in_data[532]};
    
    wire lut_637_out = lut_637_table[lut_637_select];
    
    generate
    if ( USE_REG ) begin : ff_637
        reg   lut_637_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_637_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_637_ff <= lut_637_out;
            end
        end
        
        assign out_data[637] = lut_637_ff;
    end
    else begin : no_ff_637
        assign out_data[637] = lut_637_out;
    end
    endgenerate
    
    
    
    // LUT : 638
    wire [15:0] lut_638_table = 16'b1000000011000000;
    wire [3:0] lut_638_select = {
                             in_data[550],
                             in_data[407],
                             in_data[387],
                             in_data[90]};
    
    wire lut_638_out = lut_638_table[lut_638_select];
    
    generate
    if ( USE_REG ) begin : ff_638
        reg   lut_638_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_638_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_638_ff <= lut_638_out;
            end
        end
        
        assign out_data[638] = lut_638_ff;
    end
    else begin : no_ff_638
        assign out_data[638] = lut_638_out;
    end
    endgenerate
    
    
    
    // LUT : 639
    wire [15:0] lut_639_table = 16'b0111000001110111;
    wire [3:0] lut_639_select = {
                             in_data[258],
                             in_data[399],
                             in_data[346],
                             in_data[262]};
    
    wire lut_639_out = lut_639_table[lut_639_select];
    
    generate
    if ( USE_REG ) begin : ff_639
        reg   lut_639_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_639_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_639_ff <= lut_639_out;
            end
        end
        
        assign out_data[639] = lut_639_ff;
    end
    else begin : no_ff_639
        assign out_data[639] = lut_639_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub6
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        639:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [        159:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub6_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub6_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub6_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [639:0]  in_data,
            output wire [159:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b0000000011110011;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b0100000011011101;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b0011111100000010;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b0101010011111111;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b0001011100000101;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1111101010000000;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b0000000000100011;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1111110011101000;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b0011000100010001;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b1101010011011101;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b0001011101111111;
    wire [3:0] lut_10_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b1111010100010000;
    wire [3:0] lut_11_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b0010000010110000;
    wire [3:0] lut_12_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b1100010011011100;
    wire [3:0] lut_13_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b0011111100100011;
    wire [3:0] lut_14_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b1000111000001000;
    wire [3:0] lut_15_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b1110100011101010;
    wire [3:0] lut_16_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b1101111101001101;
    wire [3:0] lut_17_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0000011101011111;
    wire [3:0] lut_18_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b0011000100010000;
    wire [3:0] lut_19_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b0100110100001100;
    wire [3:0] lut_20_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b1111111101011111;
    wire [3:0] lut_21_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b0000011100000111;
    wire [3:0] lut_22_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0000000001001100;
    wire [3:0] lut_23_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1110101011111110;
    wire [3:0] lut_24_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0111111100010111;
    wire [3:0] lut_25_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b0010101111111111;
    wire [3:0] lut_26_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1101010001000000;
    wire [3:0] lut_27_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b1111111110001110;
    wire [3:0] lut_28_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b0000001000001011;
    wire [3:0] lut_29_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b1100110100000100;
    wire [3:0] lut_30_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b1100000011001000;
    wire [3:0] lut_31_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b0111111100111111;
    wire [3:0] lut_32_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b0000110010001110;
    wire [3:0] lut_33_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1101010101010000;
    wire [3:0] lut_34_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1110110010001000;
    wire [3:0] lut_35_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b0000010111011111;
    wire [3:0] lut_36_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0000000010100000;
    wire [3:0] lut_37_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b1000000011101100;
    wire [3:0] lut_38_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b1111110111110101;
    wire [3:0] lut_39_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
    
    // LUT : 40
    wire [15:0] lut_40_table = 16'b0101111101111111;
    wire [3:0] lut_40_select = {
                             in_data[163],
                             in_data[162],
                             in_data[161],
                             in_data[160]};
    
    wire lut_40_out = lut_40_table[lut_40_select];
    
    generate
    if ( USE_REG ) begin : ff_40
        reg   lut_40_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_40_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_40_ff <= lut_40_out;
            end
        end
        
        assign out_data[40] = lut_40_ff;
    end
    else begin : no_ff_40
        assign out_data[40] = lut_40_out;
    end
    endgenerate
    
    
    
    // LUT : 41
    wire [15:0] lut_41_table = 16'b0011101100101011;
    wire [3:0] lut_41_select = {
                             in_data[167],
                             in_data[166],
                             in_data[165],
                             in_data[164]};
    
    wire lut_41_out = lut_41_table[lut_41_select];
    
    generate
    if ( USE_REG ) begin : ff_41
        reg   lut_41_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_41_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_41_ff <= lut_41_out;
            end
        end
        
        assign out_data[41] = lut_41_ff;
    end
    else begin : no_ff_41
        assign out_data[41] = lut_41_out;
    end
    endgenerate
    
    
    
    // LUT : 42
    wire [15:0] lut_42_table = 16'b1111101110110011;
    wire [3:0] lut_42_select = {
                             in_data[171],
                             in_data[170],
                             in_data[169],
                             in_data[168]};
    
    wire lut_42_out = lut_42_table[lut_42_select];
    
    generate
    if ( USE_REG ) begin : ff_42
        reg   lut_42_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_42_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_42_ff <= lut_42_out;
            end
        end
        
        assign out_data[42] = lut_42_ff;
    end
    else begin : no_ff_42
        assign out_data[42] = lut_42_out;
    end
    endgenerate
    
    
    
    // LUT : 43
    wire [15:0] lut_43_table = 16'b0111000100010000;
    wire [3:0] lut_43_select = {
                             in_data[175],
                             in_data[174],
                             in_data[173],
                             in_data[172]};
    
    wire lut_43_out = lut_43_table[lut_43_select];
    
    generate
    if ( USE_REG ) begin : ff_43
        reg   lut_43_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_43_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_43_ff <= lut_43_out;
            end
        end
        
        assign out_data[43] = lut_43_ff;
    end
    else begin : no_ff_43
        assign out_data[43] = lut_43_out;
    end
    endgenerate
    
    
    
    // LUT : 44
    wire [15:0] lut_44_table = 16'b0010001000000011;
    wire [3:0] lut_44_select = {
                             in_data[179],
                             in_data[178],
                             in_data[177],
                             in_data[176]};
    
    wire lut_44_out = lut_44_table[lut_44_select];
    
    generate
    if ( USE_REG ) begin : ff_44
        reg   lut_44_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_44_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_44_ff <= lut_44_out;
            end
        end
        
        assign out_data[44] = lut_44_ff;
    end
    else begin : no_ff_44
        assign out_data[44] = lut_44_out;
    end
    endgenerate
    
    
    
    // LUT : 45
    wire [15:0] lut_45_table = 16'b1111111110110010;
    wire [3:0] lut_45_select = {
                             in_data[183],
                             in_data[182],
                             in_data[181],
                             in_data[180]};
    
    wire lut_45_out = lut_45_table[lut_45_select];
    
    generate
    if ( USE_REG ) begin : ff_45
        reg   lut_45_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_45_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_45_ff <= lut_45_out;
            end
        end
        
        assign out_data[45] = lut_45_ff;
    end
    else begin : no_ff_45
        assign out_data[45] = lut_45_out;
    end
    endgenerate
    
    
    
    // LUT : 46
    wire [15:0] lut_46_table = 16'b1100010011011101;
    wire [3:0] lut_46_select = {
                             in_data[187],
                             in_data[186],
                             in_data[185],
                             in_data[184]};
    
    wire lut_46_out = lut_46_table[lut_46_select];
    
    generate
    if ( USE_REG ) begin : ff_46
        reg   lut_46_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_46_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_46_ff <= lut_46_out;
            end
        end
        
        assign out_data[46] = lut_46_ff;
    end
    else begin : no_ff_46
        assign out_data[46] = lut_46_out;
    end
    endgenerate
    
    
    
    // LUT : 47
    wire [15:0] lut_47_table = 16'b1101111111001010;
    wire [3:0] lut_47_select = {
                             in_data[191],
                             in_data[190],
                             in_data[189],
                             in_data[188]};
    
    wire lut_47_out = lut_47_table[lut_47_select];
    
    generate
    if ( USE_REG ) begin : ff_47
        reg   lut_47_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_47_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_47_ff <= lut_47_out;
            end
        end
        
        assign out_data[47] = lut_47_ff;
    end
    else begin : no_ff_47
        assign out_data[47] = lut_47_out;
    end
    endgenerate
    
    
    
    // LUT : 48
    wire [15:0] lut_48_table = 16'b0000101010101111;
    wire [3:0] lut_48_select = {
                             in_data[195],
                             in_data[194],
                             in_data[193],
                             in_data[192]};
    
    wire lut_48_out = lut_48_table[lut_48_select];
    
    generate
    if ( USE_REG ) begin : ff_48
        reg   lut_48_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_48_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_48_ff <= lut_48_out;
            end
        end
        
        assign out_data[48] = lut_48_ff;
    end
    else begin : no_ff_48
        assign out_data[48] = lut_48_out;
    end
    endgenerate
    
    
    
    // LUT : 49
    wire [15:0] lut_49_table = 16'b1111110111010100;
    wire [3:0] lut_49_select = {
                             in_data[199],
                             in_data[198],
                             in_data[197],
                             in_data[196]};
    
    wire lut_49_out = lut_49_table[lut_49_select];
    
    generate
    if ( USE_REG ) begin : ff_49
        reg   lut_49_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_49_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_49_ff <= lut_49_out;
            end
        end
        
        assign out_data[49] = lut_49_ff;
    end
    else begin : no_ff_49
        assign out_data[49] = lut_49_out;
    end
    endgenerate
    
    
    
    // LUT : 50
    wire [15:0] lut_50_table = 16'b0010000000100010;
    wire [3:0] lut_50_select = {
                             in_data[203],
                             in_data[202],
                             in_data[201],
                             in_data[200]};
    
    wire lut_50_out = lut_50_table[lut_50_select];
    
    generate
    if ( USE_REG ) begin : ff_50
        reg   lut_50_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_50_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_50_ff <= lut_50_out;
            end
        end
        
        assign out_data[50] = lut_50_ff;
    end
    else begin : no_ff_50
        assign out_data[50] = lut_50_out;
    end
    endgenerate
    
    
    
    // LUT : 51
    wire [15:0] lut_51_table = 16'b1111111100101111;
    wire [3:0] lut_51_select = {
                             in_data[207],
                             in_data[206],
                             in_data[205],
                             in_data[204]};
    
    wire lut_51_out = lut_51_table[lut_51_select];
    
    generate
    if ( USE_REG ) begin : ff_51
        reg   lut_51_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_51_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_51_ff <= lut_51_out;
            end
        end
        
        assign out_data[51] = lut_51_ff;
    end
    else begin : no_ff_51
        assign out_data[51] = lut_51_out;
    end
    endgenerate
    
    
    
    // LUT : 52
    wire [15:0] lut_52_table = 16'b1111111011101010;
    wire [3:0] lut_52_select = {
                             in_data[211],
                             in_data[210],
                             in_data[209],
                             in_data[208]};
    
    wire lut_52_out = lut_52_table[lut_52_select];
    
    generate
    if ( USE_REG ) begin : ff_52
        reg   lut_52_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_52_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_52_ff <= lut_52_out;
            end
        end
        
        assign out_data[52] = lut_52_ff;
    end
    else begin : no_ff_52
        assign out_data[52] = lut_52_out;
    end
    endgenerate
    
    
    
    // LUT : 53
    wire [15:0] lut_53_table = 16'b1101110111000000;
    wire [3:0] lut_53_select = {
                             in_data[215],
                             in_data[214],
                             in_data[213],
                             in_data[212]};
    
    wire lut_53_out = lut_53_table[lut_53_select];
    
    generate
    if ( USE_REG ) begin : ff_53
        reg   lut_53_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_53_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_53_ff <= lut_53_out;
            end
        end
        
        assign out_data[53] = lut_53_ff;
    end
    else begin : no_ff_53
        assign out_data[53] = lut_53_out;
    end
    endgenerate
    
    
    
    // LUT : 54
    wire [15:0] lut_54_table = 16'b1111110111000100;
    wire [3:0] lut_54_select = {
                             in_data[219],
                             in_data[218],
                             in_data[217],
                             in_data[216]};
    
    wire lut_54_out = lut_54_table[lut_54_select];
    
    generate
    if ( USE_REG ) begin : ff_54
        reg   lut_54_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_54_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_54_ff <= lut_54_out;
            end
        end
        
        assign out_data[54] = lut_54_ff;
    end
    else begin : no_ff_54
        assign out_data[54] = lut_54_out;
    end
    endgenerate
    
    
    
    // LUT : 55
    wire [15:0] lut_55_table = 16'b1111111111011100;
    wire [3:0] lut_55_select = {
                             in_data[223],
                             in_data[222],
                             in_data[221],
                             in_data[220]};
    
    wire lut_55_out = lut_55_table[lut_55_select];
    
    generate
    if ( USE_REG ) begin : ff_55
        reg   lut_55_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_55_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_55_ff <= lut_55_out;
            end
        end
        
        assign out_data[55] = lut_55_ff;
    end
    else begin : no_ff_55
        assign out_data[55] = lut_55_out;
    end
    endgenerate
    
    
    
    // LUT : 56
    wire [15:0] lut_56_table = 16'b0010001100000000;
    wire [3:0] lut_56_select = {
                             in_data[227],
                             in_data[226],
                             in_data[225],
                             in_data[224]};
    
    wire lut_56_out = lut_56_table[lut_56_select];
    
    generate
    if ( USE_REG ) begin : ff_56
        reg   lut_56_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_56_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_56_ff <= lut_56_out;
            end
        end
        
        assign out_data[56] = lut_56_ff;
    end
    else begin : no_ff_56
        assign out_data[56] = lut_56_out;
    end
    endgenerate
    
    
    
    // LUT : 57
    wire [15:0] lut_57_table = 16'b1100110110001100;
    wire [3:0] lut_57_select = {
                             in_data[231],
                             in_data[230],
                             in_data[229],
                             in_data[228]};
    
    wire lut_57_out = lut_57_table[lut_57_select];
    
    generate
    if ( USE_REG ) begin : ff_57
        reg   lut_57_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_57_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_57_ff <= lut_57_out;
            end
        end
        
        assign out_data[57] = lut_57_ff;
    end
    else begin : no_ff_57
        assign out_data[57] = lut_57_out;
    end
    endgenerate
    
    
    
    // LUT : 58
    wire [15:0] lut_58_table = 16'b0101111100000011;
    wire [3:0] lut_58_select = {
                             in_data[235],
                             in_data[234],
                             in_data[233],
                             in_data[232]};
    
    wire lut_58_out = lut_58_table[lut_58_select];
    
    generate
    if ( USE_REG ) begin : ff_58
        reg   lut_58_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_58_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_58_ff <= lut_58_out;
            end
        end
        
        assign out_data[58] = lut_58_ff;
    end
    else begin : no_ff_58
        assign out_data[58] = lut_58_out;
    end
    endgenerate
    
    
    
    // LUT : 59
    wire [15:0] lut_59_table = 16'b0000000000100011;
    wire [3:0] lut_59_select = {
                             in_data[239],
                             in_data[238],
                             in_data[237],
                             in_data[236]};
    
    wire lut_59_out = lut_59_table[lut_59_select];
    
    generate
    if ( USE_REG ) begin : ff_59
        reg   lut_59_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_59_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_59_ff <= lut_59_out;
            end
        end
        
        assign out_data[59] = lut_59_ff;
    end
    else begin : no_ff_59
        assign out_data[59] = lut_59_out;
    end
    endgenerate
    
    
    
    // LUT : 60
    wire [15:0] lut_60_table = 16'b1110111111001000;
    wire [3:0] lut_60_select = {
                             in_data[243],
                             in_data[242],
                             in_data[241],
                             in_data[240]};
    
    wire lut_60_out = lut_60_table[lut_60_select];
    
    generate
    if ( USE_REG ) begin : ff_60
        reg   lut_60_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_60_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_60_ff <= lut_60_out;
            end
        end
        
        assign out_data[60] = lut_60_ff;
    end
    else begin : no_ff_60
        assign out_data[60] = lut_60_out;
    end
    endgenerate
    
    
    
    // LUT : 61
    wire [15:0] lut_61_table = 16'b1010001010110000;
    wire [3:0] lut_61_select = {
                             in_data[247],
                             in_data[246],
                             in_data[245],
                             in_data[244]};
    
    wire lut_61_out = lut_61_table[lut_61_select];
    
    generate
    if ( USE_REG ) begin : ff_61
        reg   lut_61_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_61_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_61_ff <= lut_61_out;
            end
        end
        
        assign out_data[61] = lut_61_ff;
    end
    else begin : no_ff_61
        assign out_data[61] = lut_61_out;
    end
    endgenerate
    
    
    
    // LUT : 62
    wire [15:0] lut_62_table = 16'b0100110101001101;
    wire [3:0] lut_62_select = {
                             in_data[251],
                             in_data[250],
                             in_data[249],
                             in_data[248]};
    
    wire lut_62_out = lut_62_table[lut_62_select];
    
    generate
    if ( USE_REG ) begin : ff_62
        reg   lut_62_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_62_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_62_ff <= lut_62_out;
            end
        end
        
        assign out_data[62] = lut_62_ff;
    end
    else begin : no_ff_62
        assign out_data[62] = lut_62_out;
    end
    endgenerate
    
    
    
    // LUT : 63
    wire [15:0] lut_63_table = 16'b1111111111110000;
    wire [3:0] lut_63_select = {
                             in_data[255],
                             in_data[254],
                             in_data[253],
                             in_data[252]};
    
    wire lut_63_out = lut_63_table[lut_63_select];
    
    generate
    if ( USE_REG ) begin : ff_63
        reg   lut_63_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_63_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_63_ff <= lut_63_out;
            end
        end
        
        assign out_data[63] = lut_63_ff;
    end
    else begin : no_ff_63
        assign out_data[63] = lut_63_out;
    end
    endgenerate
    
    
    
    // LUT : 64
    wire [15:0] lut_64_table = 16'b1011001010110010;
    wire [3:0] lut_64_select = {
                             in_data[259],
                             in_data[258],
                             in_data[257],
                             in_data[256]};
    
    wire lut_64_out = lut_64_table[lut_64_select];
    
    generate
    if ( USE_REG ) begin : ff_64
        reg   lut_64_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_64_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_64_ff <= lut_64_out;
            end
        end
        
        assign out_data[64] = lut_64_ff;
    end
    else begin : no_ff_64
        assign out_data[64] = lut_64_out;
    end
    endgenerate
    
    
    
    // LUT : 65
    wire [15:0] lut_65_table = 16'b0010101111111111;
    wire [3:0] lut_65_select = {
                             in_data[263],
                             in_data[262],
                             in_data[261],
                             in_data[260]};
    
    wire lut_65_out = lut_65_table[lut_65_select];
    
    generate
    if ( USE_REG ) begin : ff_65
        reg   lut_65_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_65_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_65_ff <= lut_65_out;
            end
        end
        
        assign out_data[65] = lut_65_ff;
    end
    else begin : no_ff_65
        assign out_data[65] = lut_65_out;
    end
    endgenerate
    
    
    
    // LUT : 66
    wire [15:0] lut_66_table = 16'b1010001000000000;
    wire [3:0] lut_66_select = {
                             in_data[267],
                             in_data[266],
                             in_data[265],
                             in_data[264]};
    
    wire lut_66_out = lut_66_table[lut_66_select];
    
    generate
    if ( USE_REG ) begin : ff_66
        reg   lut_66_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_66_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_66_ff <= lut_66_out;
            end
        end
        
        assign out_data[66] = lut_66_ff;
    end
    else begin : no_ff_66
        assign out_data[66] = lut_66_out;
    end
    endgenerate
    
    
    
    // LUT : 67
    wire [15:0] lut_67_table = 16'b1010100010000000;
    wire [3:0] lut_67_select = {
                             in_data[271],
                             in_data[270],
                             in_data[269],
                             in_data[268]};
    
    wire lut_67_out = lut_67_table[lut_67_select];
    
    generate
    if ( USE_REG ) begin : ff_67
        reg   lut_67_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_67_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_67_ff <= lut_67_out;
            end
        end
        
        assign out_data[67] = lut_67_ff;
    end
    else begin : no_ff_67
        assign out_data[67] = lut_67_out;
    end
    endgenerate
    
    
    
    // LUT : 68
    wire [15:0] lut_68_table = 16'b0100000011111101;
    wire [3:0] lut_68_select = {
                             in_data[275],
                             in_data[274],
                             in_data[273],
                             in_data[272]};
    
    wire lut_68_out = lut_68_table[lut_68_select];
    
    generate
    if ( USE_REG ) begin : ff_68
        reg   lut_68_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_68_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_68_ff <= lut_68_out;
            end
        end
        
        assign out_data[68] = lut_68_ff;
    end
    else begin : no_ff_68
        assign out_data[68] = lut_68_out;
    end
    endgenerate
    
    
    
    // LUT : 69
    wire [15:0] lut_69_table = 16'b0100110101001101;
    wire [3:0] lut_69_select = {
                             in_data[279],
                             in_data[278],
                             in_data[277],
                             in_data[276]};
    
    wire lut_69_out = lut_69_table[lut_69_select];
    
    generate
    if ( USE_REG ) begin : ff_69
        reg   lut_69_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_69_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_69_ff <= lut_69_out;
            end
        end
        
        assign out_data[69] = lut_69_ff;
    end
    else begin : no_ff_69
        assign out_data[69] = lut_69_out;
    end
    endgenerate
    
    
    
    // LUT : 70
    wire [15:0] lut_70_table = 16'b1011001000100000;
    wire [3:0] lut_70_select = {
                             in_data[283],
                             in_data[282],
                             in_data[281],
                             in_data[280]};
    
    wire lut_70_out = lut_70_table[lut_70_select];
    
    generate
    if ( USE_REG ) begin : ff_70
        reg   lut_70_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_70_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_70_ff <= lut_70_out;
            end
        end
        
        assign out_data[70] = lut_70_ff;
    end
    else begin : no_ff_70
        assign out_data[70] = lut_70_out;
    end
    endgenerate
    
    
    
    // LUT : 71
    wire [15:0] lut_71_table = 16'b0000101000001000;
    wire [3:0] lut_71_select = {
                             in_data[287],
                             in_data[286],
                             in_data[285],
                             in_data[284]};
    
    wire lut_71_out = lut_71_table[lut_71_select];
    
    generate
    if ( USE_REG ) begin : ff_71
        reg   lut_71_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_71_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_71_ff <= lut_71_out;
            end
        end
        
        assign out_data[71] = lut_71_ff;
    end
    else begin : no_ff_71
        assign out_data[71] = lut_71_out;
    end
    endgenerate
    
    
    
    // LUT : 72
    wire [15:0] lut_72_table = 16'b1111110111010101;
    wire [3:0] lut_72_select = {
                             in_data[291],
                             in_data[290],
                             in_data[289],
                             in_data[288]};
    
    wire lut_72_out = lut_72_table[lut_72_select];
    
    generate
    if ( USE_REG ) begin : ff_72
        reg   lut_72_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_72_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_72_ff <= lut_72_out;
            end
        end
        
        assign out_data[72] = lut_72_ff;
    end
    else begin : no_ff_72
        assign out_data[72] = lut_72_out;
    end
    endgenerate
    
    
    
    // LUT : 73
    wire [15:0] lut_73_table = 16'b1111111100101111;
    wire [3:0] lut_73_select = {
                             in_data[295],
                             in_data[294],
                             in_data[293],
                             in_data[292]};
    
    wire lut_73_out = lut_73_table[lut_73_select];
    
    generate
    if ( USE_REG ) begin : ff_73
        reg   lut_73_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_73_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_73_ff <= lut_73_out;
            end
        end
        
        assign out_data[73] = lut_73_ff;
    end
    else begin : no_ff_73
        assign out_data[73] = lut_73_out;
    end
    endgenerate
    
    
    
    // LUT : 74
    wire [15:0] lut_74_table = 16'b0000000100010011;
    wire [3:0] lut_74_select = {
                             in_data[299],
                             in_data[298],
                             in_data[297],
                             in_data[296]};
    
    wire lut_74_out = lut_74_table[lut_74_select];
    
    generate
    if ( USE_REG ) begin : ff_74
        reg   lut_74_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_74_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_74_ff <= lut_74_out;
            end
        end
        
        assign out_data[74] = lut_74_ff;
    end
    else begin : no_ff_74
        assign out_data[74] = lut_74_out;
    end
    endgenerate
    
    
    
    // LUT : 75
    wire [15:0] lut_75_table = 16'b1000100000001010;
    wire [3:0] lut_75_select = {
                             in_data[303],
                             in_data[302],
                             in_data[301],
                             in_data[300]};
    
    wire lut_75_out = lut_75_table[lut_75_select];
    
    generate
    if ( USE_REG ) begin : ff_75
        reg   lut_75_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_75_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_75_ff <= lut_75_out;
            end
        end
        
        assign out_data[75] = lut_75_ff;
    end
    else begin : no_ff_75
        assign out_data[75] = lut_75_out;
    end
    endgenerate
    
    
    
    // LUT : 76
    wire [15:0] lut_76_table = 16'b0111010101010001;
    wire [3:0] lut_76_select = {
                             in_data[307],
                             in_data[306],
                             in_data[305],
                             in_data[304]};
    
    wire lut_76_out = lut_76_table[lut_76_select];
    
    generate
    if ( USE_REG ) begin : ff_76
        reg   lut_76_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_76_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_76_ff <= lut_76_out;
            end
        end
        
        assign out_data[76] = lut_76_ff;
    end
    else begin : no_ff_76
        assign out_data[76] = lut_76_out;
    end
    endgenerate
    
    
    
    // LUT : 77
    wire [15:0] lut_77_table = 16'b1000000011101000;
    wire [3:0] lut_77_select = {
                             in_data[311],
                             in_data[310],
                             in_data[309],
                             in_data[308]};
    
    wire lut_77_out = lut_77_table[lut_77_select];
    
    generate
    if ( USE_REG ) begin : ff_77
        reg   lut_77_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_77_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_77_ff <= lut_77_out;
            end
        end
        
        assign out_data[77] = lut_77_ff;
    end
    else begin : no_ff_77
        assign out_data[77] = lut_77_out;
    end
    endgenerate
    
    
    
    // LUT : 78
    wire [15:0] lut_78_table = 16'b0000000001110001;
    wire [3:0] lut_78_select = {
                             in_data[315],
                             in_data[314],
                             in_data[313],
                             in_data[312]};
    
    wire lut_78_out = lut_78_table[lut_78_select];
    
    generate
    if ( USE_REG ) begin : ff_78
        reg   lut_78_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_78_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_78_ff <= lut_78_out;
            end
        end
        
        assign out_data[78] = lut_78_ff;
    end
    else begin : no_ff_78
        assign out_data[78] = lut_78_out;
    end
    endgenerate
    
    
    
    // LUT : 79
    wire [15:0] lut_79_table = 16'b0000110100000101;
    wire [3:0] lut_79_select = {
                             in_data[319],
                             in_data[318],
                             in_data[317],
                             in_data[316]};
    
    wire lut_79_out = lut_79_table[lut_79_select];
    
    generate
    if ( USE_REG ) begin : ff_79
        reg   lut_79_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_79_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_79_ff <= lut_79_out;
            end
        end
        
        assign out_data[79] = lut_79_ff;
    end
    else begin : no_ff_79
        assign out_data[79] = lut_79_out;
    end
    endgenerate
    
    
    
    // LUT : 80
    wire [15:0] lut_80_table = 16'b1110101010101000;
    wire [3:0] lut_80_select = {
                             in_data[323],
                             in_data[322],
                             in_data[321],
                             in_data[320]};
    
    wire lut_80_out = lut_80_table[lut_80_select];
    
    generate
    if ( USE_REG ) begin : ff_80
        reg   lut_80_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_80_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_80_ff <= lut_80_out;
            end
        end
        
        assign out_data[80] = lut_80_ff;
    end
    else begin : no_ff_80
        assign out_data[80] = lut_80_out;
    end
    endgenerate
    
    
    
    // LUT : 81
    wire [15:0] lut_81_table = 16'b0111111100010101;
    wire [3:0] lut_81_select = {
                             in_data[327],
                             in_data[326],
                             in_data[325],
                             in_data[324]};
    
    wire lut_81_out = lut_81_table[lut_81_select];
    
    generate
    if ( USE_REG ) begin : ff_81
        reg   lut_81_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_81_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_81_ff <= lut_81_out;
            end
        end
        
        assign out_data[81] = lut_81_ff;
    end
    else begin : no_ff_81
        assign out_data[81] = lut_81_out;
    end
    endgenerate
    
    
    
    // LUT : 82
    wire [15:0] lut_82_table = 16'b1111101110110010;
    wire [3:0] lut_82_select = {
                             in_data[331],
                             in_data[330],
                             in_data[329],
                             in_data[328]};
    
    wire lut_82_out = lut_82_table[lut_82_select];
    
    generate
    if ( USE_REG ) begin : ff_82
        reg   lut_82_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_82_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_82_ff <= lut_82_out;
            end
        end
        
        assign out_data[82] = lut_82_ff;
    end
    else begin : no_ff_82
        assign out_data[82] = lut_82_out;
    end
    endgenerate
    
    
    
    // LUT : 83
    wire [15:0] lut_83_table = 16'b0000110101001101;
    wire [3:0] lut_83_select = {
                             in_data[335],
                             in_data[334],
                             in_data[333],
                             in_data[332]};
    
    wire lut_83_out = lut_83_table[lut_83_select];
    
    generate
    if ( USE_REG ) begin : ff_83
        reg   lut_83_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_83_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_83_ff <= lut_83_out;
            end
        end
        
        assign out_data[83] = lut_83_ff;
    end
    else begin : no_ff_83
        assign out_data[83] = lut_83_out;
    end
    endgenerate
    
    
    
    // LUT : 84
    wire [15:0] lut_84_table = 16'b1111001100010000;
    wire [3:0] lut_84_select = {
                             in_data[339],
                             in_data[338],
                             in_data[337],
                             in_data[336]};
    
    wire lut_84_out = lut_84_table[lut_84_select];
    
    generate
    if ( USE_REG ) begin : ff_84
        reg   lut_84_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_84_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_84_ff <= lut_84_out;
            end
        end
        
        assign out_data[84] = lut_84_ff;
    end
    else begin : no_ff_84
        assign out_data[84] = lut_84_out;
    end
    endgenerate
    
    
    
    // LUT : 85
    wire [15:0] lut_85_table = 16'b1011111100001011;
    wire [3:0] lut_85_select = {
                             in_data[343],
                             in_data[342],
                             in_data[341],
                             in_data[340]};
    
    wire lut_85_out = lut_85_table[lut_85_select];
    
    generate
    if ( USE_REG ) begin : ff_85
        reg   lut_85_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_85_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_85_ff <= lut_85_out;
            end
        end
        
        assign out_data[85] = lut_85_ff;
    end
    else begin : no_ff_85
        assign out_data[85] = lut_85_out;
    end
    endgenerate
    
    
    
    // LUT : 86
    wire [15:0] lut_86_table = 16'b0001101101111111;
    wire [3:0] lut_86_select = {
                             in_data[347],
                             in_data[346],
                             in_data[345],
                             in_data[344]};
    
    wire lut_86_out = lut_86_table[lut_86_select];
    
    generate
    if ( USE_REG ) begin : ff_86
        reg   lut_86_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_86_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_86_ff <= lut_86_out;
            end
        end
        
        assign out_data[86] = lut_86_ff;
    end
    else begin : no_ff_86
        assign out_data[86] = lut_86_out;
    end
    endgenerate
    
    
    
    // LUT : 87
    wire [15:0] lut_87_table = 16'b1000110011101111;
    wire [3:0] lut_87_select = {
                             in_data[351],
                             in_data[350],
                             in_data[349],
                             in_data[348]};
    
    wire lut_87_out = lut_87_table[lut_87_select];
    
    generate
    if ( USE_REG ) begin : ff_87
        reg   lut_87_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_87_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_87_ff <= lut_87_out;
            end
        end
        
        assign out_data[87] = lut_87_ff;
    end
    else begin : no_ff_87
        assign out_data[87] = lut_87_out;
    end
    endgenerate
    
    
    
    // LUT : 88
    wire [15:0] lut_88_table = 16'b1011101110111011;
    wire [3:0] lut_88_select = {
                             in_data[355],
                             in_data[354],
                             in_data[353],
                             in_data[352]};
    
    wire lut_88_out = lut_88_table[lut_88_select];
    
    generate
    if ( USE_REG ) begin : ff_88
        reg   lut_88_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_88_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_88_ff <= lut_88_out;
            end
        end
        
        assign out_data[88] = lut_88_ff;
    end
    else begin : no_ff_88
        assign out_data[88] = lut_88_out;
    end
    endgenerate
    
    
    
    // LUT : 89
    wire [15:0] lut_89_table = 16'b0000000001010000;
    wire [3:0] lut_89_select = {
                             in_data[359],
                             in_data[358],
                             in_data[357],
                             in_data[356]};
    
    wire lut_89_out = lut_89_table[lut_89_select];
    
    generate
    if ( USE_REG ) begin : ff_89
        reg   lut_89_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_89_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_89_ff <= lut_89_out;
            end
        end
        
        assign out_data[89] = lut_89_ff;
    end
    else begin : no_ff_89
        assign out_data[89] = lut_89_out;
    end
    endgenerate
    
    
    
    // LUT : 90
    wire [15:0] lut_90_table = 16'b0000101010101110;
    wire [3:0] lut_90_select = {
                             in_data[363],
                             in_data[362],
                             in_data[361],
                             in_data[360]};
    
    wire lut_90_out = lut_90_table[lut_90_select];
    
    generate
    if ( USE_REG ) begin : ff_90
        reg   lut_90_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_90_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_90_ff <= lut_90_out;
            end
        end
        
        assign out_data[90] = lut_90_ff;
    end
    else begin : no_ff_90
        assign out_data[90] = lut_90_out;
    end
    endgenerate
    
    
    
    // LUT : 91
    wire [15:0] lut_91_table = 16'b0010000001110000;
    wire [3:0] lut_91_select = {
                             in_data[367],
                             in_data[366],
                             in_data[365],
                             in_data[364]};
    
    wire lut_91_out = lut_91_table[lut_91_select];
    
    generate
    if ( USE_REG ) begin : ff_91
        reg   lut_91_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_91_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_91_ff <= lut_91_out;
            end
        end
        
        assign out_data[91] = lut_91_ff;
    end
    else begin : no_ff_91
        assign out_data[91] = lut_91_out;
    end
    endgenerate
    
    
    
    // LUT : 92
    wire [15:0] lut_92_table = 16'b0000100010001110;
    wire [3:0] lut_92_select = {
                             in_data[371],
                             in_data[370],
                             in_data[369],
                             in_data[368]};
    
    wire lut_92_out = lut_92_table[lut_92_select];
    
    generate
    if ( USE_REG ) begin : ff_92
        reg   lut_92_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_92_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_92_ff <= lut_92_out;
            end
        end
        
        assign out_data[92] = lut_92_ff;
    end
    else begin : no_ff_92
        assign out_data[92] = lut_92_out;
    end
    endgenerate
    
    
    
    // LUT : 93
    wire [15:0] lut_93_table = 16'b0000010001001111;
    wire [3:0] lut_93_select = {
                             in_data[375],
                             in_data[374],
                             in_data[373],
                             in_data[372]};
    
    wire lut_93_out = lut_93_table[lut_93_select];
    
    generate
    if ( USE_REG ) begin : ff_93
        reg   lut_93_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_93_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_93_ff <= lut_93_out;
            end
        end
        
        assign out_data[93] = lut_93_ff;
    end
    else begin : no_ff_93
        assign out_data[93] = lut_93_out;
    end
    endgenerate
    
    
    
    // LUT : 94
    wire [15:0] lut_94_table = 16'b1011111100111011;
    wire [3:0] lut_94_select = {
                             in_data[379],
                             in_data[378],
                             in_data[377],
                             in_data[376]};
    
    wire lut_94_out = lut_94_table[lut_94_select];
    
    generate
    if ( USE_REG ) begin : ff_94
        reg   lut_94_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_94_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_94_ff <= lut_94_out;
            end
        end
        
        assign out_data[94] = lut_94_ff;
    end
    else begin : no_ff_94
        assign out_data[94] = lut_94_out;
    end
    endgenerate
    
    
    
    // LUT : 95
    wire [15:0] lut_95_table = 16'b0101000111110101;
    wire [3:0] lut_95_select = {
                             in_data[383],
                             in_data[382],
                             in_data[381],
                             in_data[380]};
    
    wire lut_95_out = lut_95_table[lut_95_select];
    
    generate
    if ( USE_REG ) begin : ff_95
        reg   lut_95_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_95_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_95_ff <= lut_95_out;
            end
        end
        
        assign out_data[95] = lut_95_ff;
    end
    else begin : no_ff_95
        assign out_data[95] = lut_95_out;
    end
    endgenerate
    
    
    
    // LUT : 96
    wire [15:0] lut_96_table = 16'b1111101110111010;
    wire [3:0] lut_96_select = {
                             in_data[387],
                             in_data[386],
                             in_data[385],
                             in_data[384]};
    
    wire lut_96_out = lut_96_table[lut_96_select];
    
    generate
    if ( USE_REG ) begin : ff_96
        reg   lut_96_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_96_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_96_ff <= lut_96_out;
            end
        end
        
        assign out_data[96] = lut_96_ff;
    end
    else begin : no_ff_96
        assign out_data[96] = lut_96_out;
    end
    endgenerate
    
    
    
    // LUT : 97
    wire [15:0] lut_97_table = 16'b1101000001010000;
    wire [3:0] lut_97_select = {
                             in_data[391],
                             in_data[390],
                             in_data[389],
                             in_data[388]};
    
    wire lut_97_out = lut_97_table[lut_97_select];
    
    generate
    if ( USE_REG ) begin : ff_97
        reg   lut_97_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_97_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_97_ff <= lut_97_out;
            end
        end
        
        assign out_data[97] = lut_97_ff;
    end
    else begin : no_ff_97
        assign out_data[97] = lut_97_out;
    end
    endgenerate
    
    
    
    // LUT : 98
    wire [15:0] lut_98_table = 16'b1010000000000000;
    wire [3:0] lut_98_select = {
                             in_data[395],
                             in_data[394],
                             in_data[393],
                             in_data[392]};
    
    wire lut_98_out = lut_98_table[lut_98_select];
    
    generate
    if ( USE_REG ) begin : ff_98
        reg   lut_98_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_98_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_98_ff <= lut_98_out;
            end
        end
        
        assign out_data[98] = lut_98_ff;
    end
    else begin : no_ff_98
        assign out_data[98] = lut_98_out;
    end
    endgenerate
    
    
    
    // LUT : 99
    wire [15:0] lut_99_table = 16'b1000000010100000;
    wire [3:0] lut_99_select = {
                             in_data[399],
                             in_data[398],
                             in_data[397],
                             in_data[396]};
    
    wire lut_99_out = lut_99_table[lut_99_select];
    
    generate
    if ( USE_REG ) begin : ff_99
        reg   lut_99_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_99_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_99_ff <= lut_99_out;
            end
        end
        
        assign out_data[99] = lut_99_ff;
    end
    else begin : no_ff_99
        assign out_data[99] = lut_99_out;
    end
    endgenerate
    
    
    
    // LUT : 100
    wire [15:0] lut_100_table = 16'b0100110111011111;
    wire [3:0] lut_100_select = {
                             in_data[403],
                             in_data[402],
                             in_data[401],
                             in_data[400]};
    
    wire lut_100_out = lut_100_table[lut_100_select];
    
    generate
    if ( USE_REG ) begin : ff_100
        reg   lut_100_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_100_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_100_ff <= lut_100_out;
            end
        end
        
        assign out_data[100] = lut_100_ff;
    end
    else begin : no_ff_100
        assign out_data[100] = lut_100_out;
    end
    endgenerate
    
    
    
    // LUT : 101
    wire [15:0] lut_101_table = 16'b1111010011010000;
    wire [3:0] lut_101_select = {
                             in_data[407],
                             in_data[406],
                             in_data[405],
                             in_data[404]};
    
    wire lut_101_out = lut_101_table[lut_101_select];
    
    generate
    if ( USE_REG ) begin : ff_101
        reg   lut_101_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_101_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_101_ff <= lut_101_out;
            end
        end
        
        assign out_data[101] = lut_101_ff;
    end
    else begin : no_ff_101
        assign out_data[101] = lut_101_out;
    end
    endgenerate
    
    
    
    // LUT : 102
    wire [15:0] lut_102_table = 16'b0000001000101010;
    wire [3:0] lut_102_select = {
                             in_data[411],
                             in_data[410],
                             in_data[409],
                             in_data[408]};
    
    wire lut_102_out = lut_102_table[lut_102_select];
    
    generate
    if ( USE_REG ) begin : ff_102
        reg   lut_102_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_102_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_102_ff <= lut_102_out;
            end
        end
        
        assign out_data[102] = lut_102_ff;
    end
    else begin : no_ff_102
        assign out_data[102] = lut_102_out;
    end
    endgenerate
    
    
    
    // LUT : 103
    wire [15:0] lut_103_table = 16'b1010111111101111;
    wire [3:0] lut_103_select = {
                             in_data[415],
                             in_data[414],
                             in_data[413],
                             in_data[412]};
    
    wire lut_103_out = lut_103_table[lut_103_select];
    
    generate
    if ( USE_REG ) begin : ff_103
        reg   lut_103_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_103_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_103_ff <= lut_103_out;
            end
        end
        
        assign out_data[103] = lut_103_ff;
    end
    else begin : no_ff_103
        assign out_data[103] = lut_103_out;
    end
    endgenerate
    
    
    
    // LUT : 104
    wire [15:0] lut_104_table = 16'b1010000010000000;
    wire [3:0] lut_104_select = {
                             in_data[419],
                             in_data[418],
                             in_data[417],
                             in_data[416]};
    
    wire lut_104_out = lut_104_table[lut_104_select];
    
    generate
    if ( USE_REG ) begin : ff_104
        reg   lut_104_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_104_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_104_ff <= lut_104_out;
            end
        end
        
        assign out_data[104] = lut_104_ff;
    end
    else begin : no_ff_104
        assign out_data[104] = lut_104_out;
    end
    endgenerate
    
    
    
    // LUT : 105
    wire [15:0] lut_105_table = 16'b1011001000100000;
    wire [3:0] lut_105_select = {
                             in_data[423],
                             in_data[422],
                             in_data[421],
                             in_data[420]};
    
    wire lut_105_out = lut_105_table[lut_105_select];
    
    generate
    if ( USE_REG ) begin : ff_105
        reg   lut_105_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_105_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_105_ff <= lut_105_out;
            end
        end
        
        assign out_data[105] = lut_105_ff;
    end
    else begin : no_ff_105
        assign out_data[105] = lut_105_out;
    end
    endgenerate
    
    
    
    // LUT : 106
    wire [15:0] lut_106_table = 16'b0011001100100000;
    wire [3:0] lut_106_select = {
                             in_data[427],
                             in_data[426],
                             in_data[425],
                             in_data[424]};
    
    wire lut_106_out = lut_106_table[lut_106_select];
    
    generate
    if ( USE_REG ) begin : ff_106
        reg   lut_106_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_106_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_106_ff <= lut_106_out;
            end
        end
        
        assign out_data[106] = lut_106_ff;
    end
    else begin : no_ff_106
        assign out_data[106] = lut_106_out;
    end
    endgenerate
    
    
    
    // LUT : 107
    wire [15:0] lut_107_table = 16'b1111010111110101;
    wire [3:0] lut_107_select = {
                             in_data[431],
                             in_data[430],
                             in_data[429],
                             in_data[428]};
    
    wire lut_107_out = lut_107_table[lut_107_select];
    
    generate
    if ( USE_REG ) begin : ff_107
        reg   lut_107_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_107_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_107_ff <= lut_107_out;
            end
        end
        
        assign out_data[107] = lut_107_ff;
    end
    else begin : no_ff_107
        assign out_data[107] = lut_107_out;
    end
    endgenerate
    
    
    
    // LUT : 108
    wire [15:0] lut_108_table = 16'b1011111100101011;
    wire [3:0] lut_108_select = {
                             in_data[435],
                             in_data[434],
                             in_data[433],
                             in_data[432]};
    
    wire lut_108_out = lut_108_table[lut_108_select];
    
    generate
    if ( USE_REG ) begin : ff_108
        reg   lut_108_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_108_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_108_ff <= lut_108_out;
            end
        end
        
        assign out_data[108] = lut_108_ff;
    end
    else begin : no_ff_108
        assign out_data[108] = lut_108_out;
    end
    endgenerate
    
    
    
    // LUT : 109
    wire [15:0] lut_109_table = 16'b0000000100110011;
    wire [3:0] lut_109_select = {
                             in_data[439],
                             in_data[438],
                             in_data[437],
                             in_data[436]};
    
    wire lut_109_out = lut_109_table[lut_109_select];
    
    generate
    if ( USE_REG ) begin : ff_109
        reg   lut_109_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_109_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_109_ff <= lut_109_out;
            end
        end
        
        assign out_data[109] = lut_109_ff;
    end
    else begin : no_ff_109
        assign out_data[109] = lut_109_out;
    end
    endgenerate
    
    
    
    // LUT : 110
    wire [15:0] lut_110_table = 16'b0000010000001100;
    wire [3:0] lut_110_select = {
                             in_data[443],
                             in_data[442],
                             in_data[441],
                             in_data[440]};
    
    wire lut_110_out = lut_110_table[lut_110_select];
    
    generate
    if ( USE_REG ) begin : ff_110
        reg   lut_110_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_110_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_110_ff <= lut_110_out;
            end
        end
        
        assign out_data[110] = lut_110_ff;
    end
    else begin : no_ff_110
        assign out_data[110] = lut_110_out;
    end
    endgenerate
    
    
    
    // LUT : 111
    wire [15:0] lut_111_table = 16'b0000110000001111;
    wire [3:0] lut_111_select = {
                             in_data[447],
                             in_data[446],
                             in_data[445],
                             in_data[444]};
    
    wire lut_111_out = lut_111_table[lut_111_select];
    
    generate
    if ( USE_REG ) begin : ff_111
        reg   lut_111_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_111_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_111_ff <= lut_111_out;
            end
        end
        
        assign out_data[111] = lut_111_ff;
    end
    else begin : no_ff_111
        assign out_data[111] = lut_111_out;
    end
    endgenerate
    
    
    
    // LUT : 112
    wire [15:0] lut_112_table = 16'b0000001001101111;
    wire [3:0] lut_112_select = {
                             in_data[451],
                             in_data[450],
                             in_data[449],
                             in_data[448]};
    
    wire lut_112_out = lut_112_table[lut_112_select];
    
    generate
    if ( USE_REG ) begin : ff_112
        reg   lut_112_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_112_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_112_ff <= lut_112_out;
            end
        end
        
        assign out_data[112] = lut_112_ff;
    end
    else begin : no_ff_112
        assign out_data[112] = lut_112_out;
    end
    endgenerate
    
    
    
    // LUT : 113
    wire [15:0] lut_113_table = 16'b1101010001000000;
    wire [3:0] lut_113_select = {
                             in_data[455],
                             in_data[454],
                             in_data[453],
                             in_data[452]};
    
    wire lut_113_out = lut_113_table[lut_113_select];
    
    generate
    if ( USE_REG ) begin : ff_113
        reg   lut_113_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_113_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_113_ff <= lut_113_out;
            end
        end
        
        assign out_data[113] = lut_113_ff;
    end
    else begin : no_ff_113
        assign out_data[113] = lut_113_out;
    end
    endgenerate
    
    
    
    // LUT : 114
    wire [15:0] lut_114_table = 16'b1111011111110101;
    wire [3:0] lut_114_select = {
                             in_data[459],
                             in_data[458],
                             in_data[457],
                             in_data[456]};
    
    wire lut_114_out = lut_114_table[lut_114_select];
    
    generate
    if ( USE_REG ) begin : ff_114
        reg   lut_114_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_114_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_114_ff <= lut_114_out;
            end
        end
        
        assign out_data[114] = lut_114_ff;
    end
    else begin : no_ff_114
        assign out_data[114] = lut_114_out;
    end
    endgenerate
    
    
    
    // LUT : 115
    wire [15:0] lut_115_table = 16'b0001010100010111;
    wire [3:0] lut_115_select = {
                             in_data[463],
                             in_data[462],
                             in_data[461],
                             in_data[460]};
    
    wire lut_115_out = lut_115_table[lut_115_select];
    
    generate
    if ( USE_REG ) begin : ff_115
        reg   lut_115_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_115_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_115_ff <= lut_115_out;
            end
        end
        
        assign out_data[115] = lut_115_ff;
    end
    else begin : no_ff_115
        assign out_data[115] = lut_115_out;
    end
    endgenerate
    
    
    
    // LUT : 116
    wire [15:0] lut_116_table = 16'b0001111100001101;
    wire [3:0] lut_116_select = {
                             in_data[467],
                             in_data[466],
                             in_data[465],
                             in_data[464]};
    
    wire lut_116_out = lut_116_table[lut_116_select];
    
    generate
    if ( USE_REG ) begin : ff_116
        reg   lut_116_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_116_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_116_ff <= lut_116_out;
            end
        end
        
        assign out_data[116] = lut_116_ff;
    end
    else begin : no_ff_116
        assign out_data[116] = lut_116_out;
    end
    endgenerate
    
    
    
    // LUT : 117
    wire [15:0] lut_117_table = 16'b0001000101111111;
    wire [3:0] lut_117_select = {
                             in_data[471],
                             in_data[470],
                             in_data[469],
                             in_data[468]};
    
    wire lut_117_out = lut_117_table[lut_117_select];
    
    generate
    if ( USE_REG ) begin : ff_117
        reg   lut_117_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_117_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_117_ff <= lut_117_out;
            end
        end
        
        assign out_data[117] = lut_117_ff;
    end
    else begin : no_ff_117
        assign out_data[117] = lut_117_out;
    end
    endgenerate
    
    
    
    // LUT : 118
    wire [15:0] lut_118_table = 16'b1111001101110011;
    wire [3:0] lut_118_select = {
                             in_data[475],
                             in_data[474],
                             in_data[473],
                             in_data[472]};
    
    wire lut_118_out = lut_118_table[lut_118_select];
    
    generate
    if ( USE_REG ) begin : ff_118
        reg   lut_118_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_118_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_118_ff <= lut_118_out;
            end
        end
        
        assign out_data[118] = lut_118_ff;
    end
    else begin : no_ff_118
        assign out_data[118] = lut_118_out;
    end
    endgenerate
    
    
    
    // LUT : 119
    wire [15:0] lut_119_table = 16'b0000000100010011;
    wire [3:0] lut_119_select = {
                             in_data[479],
                             in_data[478],
                             in_data[477],
                             in_data[476]};
    
    wire lut_119_out = lut_119_table[lut_119_select];
    
    generate
    if ( USE_REG ) begin : ff_119
        reg   lut_119_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_119_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_119_ff <= lut_119_out;
            end
        end
        
        assign out_data[119] = lut_119_ff;
    end
    else begin : no_ff_119
        assign out_data[119] = lut_119_out;
    end
    endgenerate
    
    
    
    // LUT : 120
    wire [15:0] lut_120_table = 16'b0101111101011111;
    wire [3:0] lut_120_select = {
                             in_data[483],
                             in_data[482],
                             in_data[481],
                             in_data[480]};
    
    wire lut_120_out = lut_120_table[lut_120_select];
    
    generate
    if ( USE_REG ) begin : ff_120
        reg   lut_120_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_120_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_120_ff <= lut_120_out;
            end
        end
        
        assign out_data[120] = lut_120_ff;
    end
    else begin : no_ff_120
        assign out_data[120] = lut_120_out;
    end
    endgenerate
    
    
    
    // LUT : 121
    wire [15:0] lut_121_table = 16'b1000000010100000;
    wire [3:0] lut_121_select = {
                             in_data[487],
                             in_data[486],
                             in_data[485],
                             in_data[484]};
    
    wire lut_121_out = lut_121_table[lut_121_select];
    
    generate
    if ( USE_REG ) begin : ff_121
        reg   lut_121_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_121_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_121_ff <= lut_121_out;
            end
        end
        
        assign out_data[121] = lut_121_ff;
    end
    else begin : no_ff_121
        assign out_data[121] = lut_121_out;
    end
    endgenerate
    
    
    
    // LUT : 122
    wire [15:0] lut_122_table = 16'b0010001010111011;
    wire [3:0] lut_122_select = {
                             in_data[491],
                             in_data[490],
                             in_data[489],
                             in_data[488]};
    
    wire lut_122_out = lut_122_table[lut_122_select];
    
    generate
    if ( USE_REG ) begin : ff_122
        reg   lut_122_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_122_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_122_ff <= lut_122_out;
            end
        end
        
        assign out_data[122] = lut_122_ff;
    end
    else begin : no_ff_122
        assign out_data[122] = lut_122_out;
    end
    endgenerate
    
    
    
    // LUT : 123
    wire [15:0] lut_123_table = 16'b1011111100101011;
    wire [3:0] lut_123_select = {
                             in_data[495],
                             in_data[494],
                             in_data[493],
                             in_data[492]};
    
    wire lut_123_out = lut_123_table[lut_123_select];
    
    generate
    if ( USE_REG ) begin : ff_123
        reg   lut_123_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_123_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_123_ff <= lut_123_out;
            end
        end
        
        assign out_data[123] = lut_123_ff;
    end
    else begin : no_ff_123
        assign out_data[123] = lut_123_out;
    end
    endgenerate
    
    
    
    // LUT : 124
    wire [15:0] lut_124_table = 16'b0000000000110011;
    wire [3:0] lut_124_select = {
                             in_data[499],
                             in_data[498],
                             in_data[497],
                             in_data[496]};
    
    wire lut_124_out = lut_124_table[lut_124_select];
    
    generate
    if ( USE_REG ) begin : ff_124
        reg   lut_124_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_124_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_124_ff <= lut_124_out;
            end
        end
        
        assign out_data[124] = lut_124_ff;
    end
    else begin : no_ff_124
        assign out_data[124] = lut_124_out;
    end
    endgenerate
    
    
    
    // LUT : 125
    wire [15:0] lut_125_table = 16'b0000000010001010;
    wire [3:0] lut_125_select = {
                             in_data[503],
                             in_data[502],
                             in_data[501],
                             in_data[500]};
    
    wire lut_125_out = lut_125_table[lut_125_select];
    
    generate
    if ( USE_REG ) begin : ff_125
        reg   lut_125_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_125_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_125_ff <= lut_125_out;
            end
        end
        
        assign out_data[125] = lut_125_ff;
    end
    else begin : no_ff_125
        assign out_data[125] = lut_125_out;
    end
    endgenerate
    
    
    
    // LUT : 126
    wire [15:0] lut_126_table = 16'b1000100011111111;
    wire [3:0] lut_126_select = {
                             in_data[507],
                             in_data[506],
                             in_data[505],
                             in_data[504]};
    
    wire lut_126_out = lut_126_table[lut_126_select];
    
    generate
    if ( USE_REG ) begin : ff_126
        reg   lut_126_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_126_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_126_ff <= lut_126_out;
            end
        end
        
        assign out_data[126] = lut_126_ff;
    end
    else begin : no_ff_126
        assign out_data[126] = lut_126_out;
    end
    endgenerate
    
    
    
    // LUT : 127
    wire [15:0] lut_127_table = 16'b0001011101111111;
    wire [3:0] lut_127_select = {
                             in_data[511],
                             in_data[510],
                             in_data[509],
                             in_data[508]};
    
    wire lut_127_out = lut_127_table[lut_127_select];
    
    generate
    if ( USE_REG ) begin : ff_127
        reg   lut_127_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_127_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_127_ff <= lut_127_out;
            end
        end
        
        assign out_data[127] = lut_127_ff;
    end
    else begin : no_ff_127
        assign out_data[127] = lut_127_out;
    end
    endgenerate
    
    
    
    // LUT : 128
    wire [15:0] lut_128_table = 16'b0000000001110001;
    wire [3:0] lut_128_select = {
                             in_data[515],
                             in_data[514],
                             in_data[513],
                             in_data[512]};
    
    wire lut_128_out = lut_128_table[lut_128_select];
    
    generate
    if ( USE_REG ) begin : ff_128
        reg   lut_128_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_128_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_128_ff <= lut_128_out;
            end
        end
        
        assign out_data[128] = lut_128_ff;
    end
    else begin : no_ff_128
        assign out_data[128] = lut_128_out;
    end
    endgenerate
    
    
    
    // LUT : 129
    wire [15:0] lut_129_table = 16'b1011001011111011;
    wire [3:0] lut_129_select = {
                             in_data[519],
                             in_data[518],
                             in_data[517],
                             in_data[516]};
    
    wire lut_129_out = lut_129_table[lut_129_select];
    
    generate
    if ( USE_REG ) begin : ff_129
        reg   lut_129_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_129_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_129_ff <= lut_129_out;
            end
        end
        
        assign out_data[129] = lut_129_ff;
    end
    else begin : no_ff_129
        assign out_data[129] = lut_129_out;
    end
    endgenerate
    
    
    
    // LUT : 130
    wire [15:0] lut_130_table = 16'b1111111111010100;
    wire [3:0] lut_130_select = {
                             in_data[523],
                             in_data[522],
                             in_data[521],
                             in_data[520]};
    
    wire lut_130_out = lut_130_table[lut_130_select];
    
    generate
    if ( USE_REG ) begin : ff_130
        reg   lut_130_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_130_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_130_ff <= lut_130_out;
            end
        end
        
        assign out_data[130] = lut_130_ff;
    end
    else begin : no_ff_130
        assign out_data[130] = lut_130_out;
    end
    endgenerate
    
    
    
    // LUT : 131
    wire [15:0] lut_131_table = 16'b1101010000000000;
    wire [3:0] lut_131_select = {
                             in_data[527],
                             in_data[526],
                             in_data[525],
                             in_data[524]};
    
    wire lut_131_out = lut_131_table[lut_131_select];
    
    generate
    if ( USE_REG ) begin : ff_131
        reg   lut_131_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_131_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_131_ff <= lut_131_out;
            end
        end
        
        assign out_data[131] = lut_131_ff;
    end
    else begin : no_ff_131
        assign out_data[131] = lut_131_out;
    end
    endgenerate
    
    
    
    // LUT : 132
    wire [15:0] lut_132_table = 16'b1100111100001100;
    wire [3:0] lut_132_select = {
                             in_data[531],
                             in_data[530],
                             in_data[529],
                             in_data[528]};
    
    wire lut_132_out = lut_132_table[lut_132_select];
    
    generate
    if ( USE_REG ) begin : ff_132
        reg   lut_132_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_132_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_132_ff <= lut_132_out;
            end
        end
        
        assign out_data[132] = lut_132_ff;
    end
    else begin : no_ff_132
        assign out_data[132] = lut_132_out;
    end
    endgenerate
    
    
    
    // LUT : 133
    wire [15:0] lut_133_table = 16'b0000101000000000;
    wire [3:0] lut_133_select = {
                             in_data[535],
                             in_data[534],
                             in_data[533],
                             in_data[532]};
    
    wire lut_133_out = lut_133_table[lut_133_select];
    
    generate
    if ( USE_REG ) begin : ff_133
        reg   lut_133_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_133_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_133_ff <= lut_133_out;
            end
        end
        
        assign out_data[133] = lut_133_ff;
    end
    else begin : no_ff_133
        assign out_data[133] = lut_133_out;
    end
    endgenerate
    
    
    
    // LUT : 134
    wire [15:0] lut_134_table = 16'b1111101110110010;
    wire [3:0] lut_134_select = {
                             in_data[539],
                             in_data[538],
                             in_data[537],
                             in_data[536]};
    
    wire lut_134_out = lut_134_table[lut_134_select];
    
    generate
    if ( USE_REG ) begin : ff_134
        reg   lut_134_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_134_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_134_ff <= lut_134_out;
            end
        end
        
        assign out_data[134] = lut_134_ff;
    end
    else begin : no_ff_134
        assign out_data[134] = lut_134_out;
    end
    endgenerate
    
    
    
    // LUT : 135
    wire [15:0] lut_135_table = 16'b0001000001010001;
    wire [3:0] lut_135_select = {
                             in_data[543],
                             in_data[542],
                             in_data[541],
                             in_data[540]};
    
    wire lut_135_out = lut_135_table[lut_135_select];
    
    generate
    if ( USE_REG ) begin : ff_135
        reg   lut_135_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_135_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_135_ff <= lut_135_out;
            end
        end
        
        assign out_data[135] = lut_135_ff;
    end
    else begin : no_ff_135
        assign out_data[135] = lut_135_out;
    end
    endgenerate
    
    
    
    // LUT : 136
    wire [15:0] lut_136_table = 16'b1101111101001100;
    wire [3:0] lut_136_select = {
                             in_data[547],
                             in_data[546],
                             in_data[545],
                             in_data[544]};
    
    wire lut_136_out = lut_136_table[lut_136_select];
    
    generate
    if ( USE_REG ) begin : ff_136
        reg   lut_136_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_136_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_136_ff <= lut_136_out;
            end
        end
        
        assign out_data[136] = lut_136_ff;
    end
    else begin : no_ff_136
        assign out_data[136] = lut_136_out;
    end
    endgenerate
    
    
    
    // LUT : 137
    wire [15:0] lut_137_table = 16'b0011000101110000;
    wire [3:0] lut_137_select = {
                             in_data[551],
                             in_data[550],
                             in_data[549],
                             in_data[548]};
    
    wire lut_137_out = lut_137_table[lut_137_select];
    
    generate
    if ( USE_REG ) begin : ff_137
        reg   lut_137_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_137_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_137_ff <= lut_137_out;
            end
        end
        
        assign out_data[137] = lut_137_ff;
    end
    else begin : no_ff_137
        assign out_data[137] = lut_137_out;
    end
    endgenerate
    
    
    
    // LUT : 138
    wire [15:0] lut_138_table = 16'b1000000010000000;
    wire [3:0] lut_138_select = {
                             in_data[555],
                             in_data[554],
                             in_data[553],
                             in_data[552]};
    
    wire lut_138_out = lut_138_table[lut_138_select];
    
    generate
    if ( USE_REG ) begin : ff_138
        reg   lut_138_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_138_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_138_ff <= lut_138_out;
            end
        end
        
        assign out_data[138] = lut_138_ff;
    end
    else begin : no_ff_138
        assign out_data[138] = lut_138_out;
    end
    endgenerate
    
    
    
    // LUT : 139
    wire [15:0] lut_139_table = 16'b0001011100000100;
    wire [3:0] lut_139_select = {
                             in_data[559],
                             in_data[558],
                             in_data[557],
                             in_data[556]};
    
    wire lut_139_out = lut_139_table[lut_139_select];
    
    generate
    if ( USE_REG ) begin : ff_139
        reg   lut_139_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_139_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_139_ff <= lut_139_out;
            end
        end
        
        assign out_data[139] = lut_139_ff;
    end
    else begin : no_ff_139
        assign out_data[139] = lut_139_out;
    end
    endgenerate
    
    
    
    // LUT : 140
    wire [15:0] lut_140_table = 16'b1000100010001000;
    wire [3:0] lut_140_select = {
                             in_data[563],
                             in_data[562],
                             in_data[561],
                             in_data[560]};
    
    wire lut_140_out = lut_140_table[lut_140_select];
    
    generate
    if ( USE_REG ) begin : ff_140
        reg   lut_140_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_140_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_140_ff <= lut_140_out;
            end
        end
        
        assign out_data[140] = lut_140_ff;
    end
    else begin : no_ff_140
        assign out_data[140] = lut_140_out;
    end
    endgenerate
    
    
    
    // LUT : 141
    wire [15:0] lut_141_table = 16'b0100000000000000;
    wire [3:0] lut_141_select = {
                             in_data[567],
                             in_data[566],
                             in_data[565],
                             in_data[564]};
    
    wire lut_141_out = lut_141_table[lut_141_select];
    
    generate
    if ( USE_REG ) begin : ff_141
        reg   lut_141_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_141_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_141_ff <= lut_141_out;
            end
        end
        
        assign out_data[141] = lut_141_ff;
    end
    else begin : no_ff_141
        assign out_data[141] = lut_141_out;
    end
    endgenerate
    
    
    
    // LUT : 142
    wire [15:0] lut_142_table = 16'b1110110011111110;
    wire [3:0] lut_142_select = {
                             in_data[571],
                             in_data[570],
                             in_data[569],
                             in_data[568]};
    
    wire lut_142_out = lut_142_table[lut_142_select];
    
    generate
    if ( USE_REG ) begin : ff_142
        reg   lut_142_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_142_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_142_ff <= lut_142_out;
            end
        end
        
        assign out_data[142] = lut_142_ff;
    end
    else begin : no_ff_142
        assign out_data[142] = lut_142_out;
    end
    endgenerate
    
    
    
    // LUT : 143
    wire [15:0] lut_143_table = 16'b0000001100000000;
    wire [3:0] lut_143_select = {
                             in_data[575],
                             in_data[574],
                             in_data[573],
                             in_data[572]};
    
    wire lut_143_out = lut_143_table[lut_143_select];
    
    generate
    if ( USE_REG ) begin : ff_143
        reg   lut_143_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_143_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_143_ff <= lut_143_out;
            end
        end
        
        assign out_data[143] = lut_143_ff;
    end
    else begin : no_ff_143
        assign out_data[143] = lut_143_out;
    end
    endgenerate
    
    
    
    // LUT : 144
    wire [15:0] lut_144_table = 16'b0000101010001111;
    wire [3:0] lut_144_select = {
                             in_data[579],
                             in_data[578],
                             in_data[577],
                             in_data[576]};
    
    wire lut_144_out = lut_144_table[lut_144_select];
    
    generate
    if ( USE_REG ) begin : ff_144
        reg   lut_144_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_144_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_144_ff <= lut_144_out;
            end
        end
        
        assign out_data[144] = lut_144_ff;
    end
    else begin : no_ff_144
        assign out_data[144] = lut_144_out;
    end
    endgenerate
    
    
    
    // LUT : 145
    wire [15:0] lut_145_table = 16'b0111000000000000;
    wire [3:0] lut_145_select = {
                             in_data[583],
                             in_data[582],
                             in_data[581],
                             in_data[580]};
    
    wire lut_145_out = lut_145_table[lut_145_select];
    
    generate
    if ( USE_REG ) begin : ff_145
        reg   lut_145_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_145_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_145_ff <= lut_145_out;
            end
        end
        
        assign out_data[145] = lut_145_ff;
    end
    else begin : no_ff_145
        assign out_data[145] = lut_145_out;
    end
    endgenerate
    
    
    
    // LUT : 146
    wire [15:0] lut_146_table = 16'b1011001010110010;
    wire [3:0] lut_146_select = {
                             in_data[587],
                             in_data[586],
                             in_data[585],
                             in_data[584]};
    
    wire lut_146_out = lut_146_table[lut_146_select];
    
    generate
    if ( USE_REG ) begin : ff_146
        reg   lut_146_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_146_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_146_ff <= lut_146_out;
            end
        end
        
        assign out_data[146] = lut_146_ff;
    end
    else begin : no_ff_146
        assign out_data[146] = lut_146_out;
    end
    endgenerate
    
    
    
    // LUT : 147
    wire [15:0] lut_147_table = 16'b0010001000001011;
    wire [3:0] lut_147_select = {
                             in_data[591],
                             in_data[590],
                             in_data[589],
                             in_data[588]};
    
    wire lut_147_out = lut_147_table[lut_147_select];
    
    generate
    if ( USE_REG ) begin : ff_147
        reg   lut_147_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_147_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_147_ff <= lut_147_out;
            end
        end
        
        assign out_data[147] = lut_147_ff;
    end
    else begin : no_ff_147
        assign out_data[147] = lut_147_out;
    end
    endgenerate
    
    
    
    // LUT : 148
    wire [15:0] lut_148_table = 16'b1111011101010000;
    wire [3:0] lut_148_select = {
                             in_data[595],
                             in_data[594],
                             in_data[593],
                             in_data[592]};
    
    wire lut_148_out = lut_148_table[lut_148_select];
    
    generate
    if ( USE_REG ) begin : ff_148
        reg   lut_148_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_148_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_148_ff <= lut_148_out;
            end
        end
        
        assign out_data[148] = lut_148_ff;
    end
    else begin : no_ff_148
        assign out_data[148] = lut_148_out;
    end
    endgenerate
    
    
    
    // LUT : 149
    wire [15:0] lut_149_table = 16'b1111111111101000;
    wire [3:0] lut_149_select = {
                             in_data[599],
                             in_data[598],
                             in_data[597],
                             in_data[596]};
    
    wire lut_149_out = lut_149_table[lut_149_select];
    
    generate
    if ( USE_REG ) begin : ff_149
        reg   lut_149_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_149_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_149_ff <= lut_149_out;
            end
        end
        
        assign out_data[149] = lut_149_ff;
    end
    else begin : no_ff_149
        assign out_data[149] = lut_149_out;
    end
    endgenerate
    
    
    
    // LUT : 150
    wire [15:0] lut_150_table = 16'b0000000010001000;
    wire [3:0] lut_150_select = {
                             in_data[603],
                             in_data[602],
                             in_data[601],
                             in_data[600]};
    
    wire lut_150_out = lut_150_table[lut_150_select];
    
    generate
    if ( USE_REG ) begin : ff_150
        reg   lut_150_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_150_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_150_ff <= lut_150_out;
            end
        end
        
        assign out_data[150] = lut_150_ff;
    end
    else begin : no_ff_150
        assign out_data[150] = lut_150_out;
    end
    endgenerate
    
    
    
    // LUT : 151
    wire [15:0] lut_151_table = 16'b0011101010111111;
    wire [3:0] lut_151_select = {
                             in_data[607],
                             in_data[606],
                             in_data[605],
                             in_data[604]};
    
    wire lut_151_out = lut_151_table[lut_151_select];
    
    generate
    if ( USE_REG ) begin : ff_151
        reg   lut_151_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_151_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_151_ff <= lut_151_out;
            end
        end
        
        assign out_data[151] = lut_151_ff;
    end
    else begin : no_ff_151
        assign out_data[151] = lut_151_out;
    end
    endgenerate
    
    
    
    // LUT : 152
    wire [15:0] lut_152_table = 16'b0000000000110011;
    wire [3:0] lut_152_select = {
                             in_data[611],
                             in_data[610],
                             in_data[609],
                             in_data[608]};
    
    wire lut_152_out = lut_152_table[lut_152_select];
    
    generate
    if ( USE_REG ) begin : ff_152
        reg   lut_152_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_152_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_152_ff <= lut_152_out;
            end
        end
        
        assign out_data[152] = lut_152_ff;
    end
    else begin : no_ff_152
        assign out_data[152] = lut_152_out;
    end
    endgenerate
    
    
    
    // LUT : 153
    wire [15:0] lut_153_table = 16'b1111111110110010;
    wire [3:0] lut_153_select = {
                             in_data[615],
                             in_data[614],
                             in_data[613],
                             in_data[612]};
    
    wire lut_153_out = lut_153_table[lut_153_select];
    
    generate
    if ( USE_REG ) begin : ff_153
        reg   lut_153_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_153_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_153_ff <= lut_153_out;
            end
        end
        
        assign out_data[153] = lut_153_ff;
    end
    else begin : no_ff_153
        assign out_data[153] = lut_153_out;
    end
    endgenerate
    
    
    
    // LUT : 154
    wire [15:0] lut_154_table = 16'b0111011100110111;
    wire [3:0] lut_154_select = {
                             in_data[619],
                             in_data[618],
                             in_data[617],
                             in_data[616]};
    
    wire lut_154_out = lut_154_table[lut_154_select];
    
    generate
    if ( USE_REG ) begin : ff_154
        reg   lut_154_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_154_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_154_ff <= lut_154_out;
            end
        end
        
        assign out_data[154] = lut_154_ff;
    end
    else begin : no_ff_154
        assign out_data[154] = lut_154_out;
    end
    endgenerate
    
    
    
    // LUT : 155
    wire [15:0] lut_155_table = 16'b1011000011111011;
    wire [3:0] lut_155_select = {
                             in_data[623],
                             in_data[622],
                             in_data[621],
                             in_data[620]};
    
    wire lut_155_out = lut_155_table[lut_155_select];
    
    generate
    if ( USE_REG ) begin : ff_155
        reg   lut_155_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_155_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_155_ff <= lut_155_out;
            end
        end
        
        assign out_data[155] = lut_155_ff;
    end
    else begin : no_ff_155
        assign out_data[155] = lut_155_out;
    end
    endgenerate
    
    
    
    // LUT : 156
    wire [15:0] lut_156_table = 16'b0000000101111111;
    wire [3:0] lut_156_select = {
                             in_data[627],
                             in_data[626],
                             in_data[625],
                             in_data[624]};
    
    wire lut_156_out = lut_156_table[lut_156_select];
    
    generate
    if ( USE_REG ) begin : ff_156
        reg   lut_156_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_156_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_156_ff <= lut_156_out;
            end
        end
        
        assign out_data[156] = lut_156_ff;
    end
    else begin : no_ff_156
        assign out_data[156] = lut_156_out;
    end
    endgenerate
    
    
    
    // LUT : 157
    wire [15:0] lut_157_table = 16'b1010111011101111;
    wire [3:0] lut_157_select = {
                             in_data[631],
                             in_data[630],
                             in_data[629],
                             in_data[628]};
    
    wire lut_157_out = lut_157_table[lut_157_select];
    
    generate
    if ( USE_REG ) begin : ff_157
        reg   lut_157_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_157_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_157_ff <= lut_157_out;
            end
        end
        
        assign out_data[157] = lut_157_ff;
    end
    else begin : no_ff_157
        assign out_data[157] = lut_157_out;
    end
    endgenerate
    
    
    
    // LUT : 158
    wire [15:0] lut_158_table = 16'b1011111110111011;
    wire [3:0] lut_158_select = {
                             in_data[635],
                             in_data[634],
                             in_data[633],
                             in_data[632]};
    
    wire lut_158_out = lut_158_table[lut_158_select];
    
    generate
    if ( USE_REG ) begin : ff_158
        reg   lut_158_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_158_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_158_ff <= lut_158_out;
            end
        end
        
        assign out_data[158] = lut_158_ff;
    end
    else begin : no_ff_158
        assign out_data[158] = lut_158_out;
    end
    endgenerate
    
    
    
    // LUT : 159
    wire [15:0] lut_159_table = 16'b0000001100111111;
    wire [3:0] lut_159_select = {
                             in_data[639],
                             in_data[638],
                             in_data[637],
                             in_data[636]};
    
    wire lut_159_out = lut_159_table[lut_159_select];
    
    generate
    if ( USE_REG ) begin : ff_159
        reg   lut_159_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_159_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_159_ff <= lut_159_out;
            end
        end
        
        assign out_data[159] = lut_159_ff;
    end
    else begin : no_ff_159
        assign out_data[159] = lut_159_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub7
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [        159:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [         39:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub7_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub7_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub7_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [159:0]  in_data,
            output wire [39:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1000000011101000;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b0100000011010100;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b0010101100000010;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1000111010001000;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b0001011100000001;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1011001010110000;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b0000000100010111;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1101010001000000;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1101010001000000;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b0100000011110100;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
    
    // LUT : 10
    wire [15:0] lut_10_table = 16'b0101011100010001;
    wire [3:0] lut_10_select = {
                             in_data[43],
                             in_data[42],
                             in_data[41],
                             in_data[40]};
    
    wire lut_10_out = lut_10_table[lut_10_select];
    
    generate
    if ( USE_REG ) begin : ff_10
        reg   lut_10_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_10_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_10_ff <= lut_10_out;
            end
        end
        
        assign out_data[10] = lut_10_ff;
    end
    else begin : no_ff_10
        assign out_data[10] = lut_10_out;
    end
    endgenerate
    
    
    
    // LUT : 11
    wire [15:0] lut_11_table = 16'b1011001000100000;
    wire [3:0] lut_11_select = {
                             in_data[47],
                             in_data[46],
                             in_data[45],
                             in_data[44]};
    
    wire lut_11_out = lut_11_table[lut_11_select];
    
    generate
    if ( USE_REG ) begin : ff_11
        reg   lut_11_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_11_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_11_ff <= lut_11_out;
            end
        end
        
        assign out_data[11] = lut_11_ff;
    end
    else begin : no_ff_11
        assign out_data[11] = lut_11_out;
    end
    endgenerate
    
    
    
    // LUT : 12
    wire [15:0] lut_12_table = 16'b0011000111110011;
    wire [3:0] lut_12_select = {
                             in_data[51],
                             in_data[50],
                             in_data[49],
                             in_data[48]};
    
    wire lut_12_out = lut_12_table[lut_12_select];
    
    generate
    if ( USE_REG ) begin : ff_12
        reg   lut_12_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_12_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_12_ff <= lut_12_out;
            end
        end
        
        assign out_data[12] = lut_12_ff;
    end
    else begin : no_ff_12
        assign out_data[12] = lut_12_out;
    end
    endgenerate
    
    
    
    // LUT : 13
    wire [15:0] lut_13_table = 16'b0000110001001101;
    wire [3:0] lut_13_select = {
                             in_data[55],
                             in_data[54],
                             in_data[53],
                             in_data[52]};
    
    wire lut_13_out = lut_13_table[lut_13_select];
    
    generate
    if ( USE_REG ) begin : ff_13
        reg   lut_13_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_13_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_13_ff <= lut_13_out;
            end
        end
        
        assign out_data[13] = lut_13_ff;
    end
    else begin : no_ff_13
        assign out_data[13] = lut_13_out;
    end
    endgenerate
    
    
    
    // LUT : 14
    wire [15:0] lut_14_table = 16'b1011001000100000;
    wire [3:0] lut_14_select = {
                             in_data[59],
                             in_data[58],
                             in_data[57],
                             in_data[56]};
    
    wire lut_14_out = lut_14_table[lut_14_select];
    
    generate
    if ( USE_REG ) begin : ff_14
        reg   lut_14_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_14_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_14_ff <= lut_14_out;
            end
        end
        
        assign out_data[14] = lut_14_ff;
    end
    else begin : no_ff_14
        assign out_data[14] = lut_14_out;
    end
    endgenerate
    
    
    
    // LUT : 15
    wire [15:0] lut_15_table = 16'b0100010011010100;
    wire [3:0] lut_15_select = {
                             in_data[63],
                             in_data[62],
                             in_data[61],
                             in_data[60]};
    
    wire lut_15_out = lut_15_table[lut_15_select];
    
    generate
    if ( USE_REG ) begin : ff_15
        reg   lut_15_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_15_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_15_ff <= lut_15_out;
            end
        end
        
        assign out_data[15] = lut_15_ff;
    end
    else begin : no_ff_15
        assign out_data[15] = lut_15_out;
    end
    endgenerate
    
    
    
    // LUT : 16
    wire [15:0] lut_16_table = 16'b1011001000100000;
    wire [3:0] lut_16_select = {
                             in_data[67],
                             in_data[66],
                             in_data[65],
                             in_data[64]};
    
    wire lut_16_out = lut_16_table[lut_16_select];
    
    generate
    if ( USE_REG ) begin : ff_16
        reg   lut_16_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_16_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_16_ff <= lut_16_out;
            end
        end
        
        assign out_data[16] = lut_16_ff;
    end
    else begin : no_ff_16
        assign out_data[16] = lut_16_out;
    end
    endgenerate
    
    
    
    // LUT : 17
    wire [15:0] lut_17_table = 16'b1101010001000000;
    wire [3:0] lut_17_select = {
                             in_data[71],
                             in_data[70],
                             in_data[69],
                             in_data[68]};
    
    wire lut_17_out = lut_17_table[lut_17_select];
    
    generate
    if ( USE_REG ) begin : ff_17
        reg   lut_17_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_17_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_17_ff <= lut_17_out;
            end
        end
        
        assign out_data[17] = lut_17_ff;
    end
    else begin : no_ff_17
        assign out_data[17] = lut_17_out;
    end
    endgenerate
    
    
    
    // LUT : 18
    wire [15:0] lut_18_table = 16'b0001000001110111;
    wire [3:0] lut_18_select = {
                             in_data[75],
                             in_data[74],
                             in_data[73],
                             in_data[72]};
    
    wire lut_18_out = lut_18_table[lut_18_select];
    
    generate
    if ( USE_REG ) begin : ff_18
        reg   lut_18_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_18_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_18_ff <= lut_18_out;
            end
        end
        
        assign out_data[18] = lut_18_ff;
    end
    else begin : no_ff_18
        assign out_data[18] = lut_18_out;
    end
    endgenerate
    
    
    
    // LUT : 19
    wire [15:0] lut_19_table = 16'b1101010001000000;
    wire [3:0] lut_19_select = {
                             in_data[79],
                             in_data[78],
                             in_data[77],
                             in_data[76]};
    
    wire lut_19_out = lut_19_table[lut_19_select];
    
    generate
    if ( USE_REG ) begin : ff_19
        reg   lut_19_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_19_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_19_ff <= lut_19_out;
            end
        end
        
        assign out_data[19] = lut_19_ff;
    end
    else begin : no_ff_19
        assign out_data[19] = lut_19_out;
    end
    endgenerate
    
    
    
    // LUT : 20
    wire [15:0] lut_20_table = 16'b1100110100001100;
    wire [3:0] lut_20_select = {
                             in_data[83],
                             in_data[82],
                             in_data[81],
                             in_data[80]};
    
    wire lut_20_out = lut_20_table[lut_20_select];
    
    generate
    if ( USE_REG ) begin : ff_20
        reg   lut_20_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_20_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_20_ff <= lut_20_out;
            end
        end
        
        assign out_data[20] = lut_20_ff;
    end
    else begin : no_ff_20
        assign out_data[20] = lut_20_out;
    end
    endgenerate
    
    
    
    // LUT : 21
    wire [15:0] lut_21_table = 16'b0100110100000100;
    wire [3:0] lut_21_select = {
                             in_data[87],
                             in_data[86],
                             in_data[85],
                             in_data[84]};
    
    wire lut_21_out = lut_21_table[lut_21_select];
    
    generate
    if ( USE_REG ) begin : ff_21
        reg   lut_21_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_21_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_21_ff <= lut_21_out;
            end
        end
        
        assign out_data[21] = lut_21_ff;
    end
    else begin : no_ff_21
        assign out_data[21] = lut_21_out;
    end
    endgenerate
    
    
    
    // LUT : 22
    wire [15:0] lut_22_table = 16'b0000010001011101;
    wire [3:0] lut_22_select = {
                             in_data[91],
                             in_data[90],
                             in_data[89],
                             in_data[88]};
    
    wire lut_22_out = lut_22_table[lut_22_select];
    
    generate
    if ( USE_REG ) begin : ff_22
        reg   lut_22_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_22_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_22_ff <= lut_22_out;
            end
        end
        
        assign out_data[22] = lut_22_ff;
    end
    else begin : no_ff_22
        assign out_data[22] = lut_22_out;
    end
    endgenerate
    
    
    
    // LUT : 23
    wire [15:0] lut_23_table = 16'b0000100010001110;
    wire [3:0] lut_23_select = {
                             in_data[95],
                             in_data[94],
                             in_data[93],
                             in_data[92]};
    
    wire lut_23_out = lut_23_table[lut_23_select];
    
    generate
    if ( USE_REG ) begin : ff_23
        reg   lut_23_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_23_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_23_ff <= lut_23_out;
            end
        end
        
        assign out_data[23] = lut_23_ff;
    end
    else begin : no_ff_23
        assign out_data[23] = lut_23_out;
    end
    endgenerate
    
    
    
    // LUT : 24
    wire [15:0] lut_24_table = 16'b1101110101000000;
    wire [3:0] lut_24_select = {
                             in_data[99],
                             in_data[98],
                             in_data[97],
                             in_data[96]};
    
    wire lut_24_out = lut_24_table[lut_24_select];
    
    generate
    if ( USE_REG ) begin : ff_24
        reg   lut_24_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_24_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_24_ff <= lut_24_out;
            end
        end
        
        assign out_data[24] = lut_24_ff;
    end
    else begin : no_ff_24
        assign out_data[24] = lut_24_out;
    end
    endgenerate
    
    
    
    // LUT : 25
    wire [15:0] lut_25_table = 16'b0001000001110001;
    wire [3:0] lut_25_select = {
                             in_data[103],
                             in_data[102],
                             in_data[101],
                             in_data[100]};
    
    wire lut_25_out = lut_25_table[lut_25_select];
    
    generate
    if ( USE_REG ) begin : ff_25
        reg   lut_25_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_25_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_25_ff <= lut_25_out;
            end
        end
        
        assign out_data[25] = lut_25_ff;
    end
    else begin : no_ff_25
        assign out_data[25] = lut_25_out;
    end
    endgenerate
    
    
    
    // LUT : 26
    wire [15:0] lut_26_table = 16'b1000000011101010;
    wire [3:0] lut_26_select = {
                             in_data[107],
                             in_data[106],
                             in_data[105],
                             in_data[104]};
    
    wire lut_26_out = lut_26_table[lut_26_select];
    
    generate
    if ( USE_REG ) begin : ff_26
        reg   lut_26_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_26_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_26_ff <= lut_26_out;
            end
        end
        
        assign out_data[26] = lut_26_ff;
    end
    else begin : no_ff_26
        assign out_data[26] = lut_26_out;
    end
    endgenerate
    
    
    
    // LUT : 27
    wire [15:0] lut_27_table = 16'b1110100010000000;
    wire [3:0] lut_27_select = {
                             in_data[111],
                             in_data[110],
                             in_data[109],
                             in_data[108]};
    
    wire lut_27_out = lut_27_table[lut_27_select];
    
    generate
    if ( USE_REG ) begin : ff_27
        reg   lut_27_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_27_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_27_ff <= lut_27_out;
            end
        end
        
        assign out_data[27] = lut_27_ff;
    end
    else begin : no_ff_27
        assign out_data[27] = lut_27_out;
    end
    endgenerate
    
    
    
    // LUT : 28
    wire [15:0] lut_28_table = 16'b1000111000001000;
    wire [3:0] lut_28_select = {
                             in_data[115],
                             in_data[114],
                             in_data[113],
                             in_data[112]};
    
    wire lut_28_out = lut_28_table[lut_28_select];
    
    generate
    if ( USE_REG ) begin : ff_28
        reg   lut_28_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_28_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_28_ff <= lut_28_out;
            end
        end
        
        assign out_data[28] = lut_28_ff;
    end
    else begin : no_ff_28
        assign out_data[28] = lut_28_out;
    end
    endgenerate
    
    
    
    // LUT : 29
    wire [15:0] lut_29_table = 16'b1000111000001000;
    wire [3:0] lut_29_select = {
                             in_data[119],
                             in_data[118],
                             in_data[117],
                             in_data[116]};
    
    wire lut_29_out = lut_29_table[lut_29_select];
    
    generate
    if ( USE_REG ) begin : ff_29
        reg   lut_29_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_29_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_29_ff <= lut_29_out;
            end
        end
        
        assign out_data[29] = lut_29_ff;
    end
    else begin : no_ff_29
        assign out_data[29] = lut_29_out;
    end
    endgenerate
    
    
    
    // LUT : 30
    wire [15:0] lut_30_table = 16'b0000010001001101;
    wire [3:0] lut_30_select = {
                             in_data[123],
                             in_data[122],
                             in_data[121],
                             in_data[120]};
    
    wire lut_30_out = lut_30_table[lut_30_select];
    
    generate
    if ( USE_REG ) begin : ff_30
        reg   lut_30_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_30_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_30_ff <= lut_30_out;
            end
        end
        
        assign out_data[30] = lut_30_ff;
    end
    else begin : no_ff_30
        assign out_data[30] = lut_30_out;
    end
    endgenerate
    
    
    
    // LUT : 31
    wire [15:0] lut_31_table = 16'b0000100010101110;
    wire [3:0] lut_31_select = {
                             in_data[127],
                             in_data[126],
                             in_data[125],
                             in_data[124]};
    
    wire lut_31_out = lut_31_table[lut_31_select];
    
    generate
    if ( USE_REG ) begin : ff_31
        reg   lut_31_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_31_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_31_ff <= lut_31_out;
            end
        end
        
        assign out_data[31] = lut_31_ff;
    end
    else begin : no_ff_31
        assign out_data[31] = lut_31_out;
    end
    endgenerate
    
    
    
    // LUT : 32
    wire [15:0] lut_32_table = 16'b0010101100000010;
    wire [3:0] lut_32_select = {
                             in_data[131],
                             in_data[130],
                             in_data[129],
                             in_data[128]};
    
    wire lut_32_out = lut_32_table[lut_32_select];
    
    generate
    if ( USE_REG ) begin : ff_32
        reg   lut_32_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_32_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_32_ff <= lut_32_out;
            end
        end
        
        assign out_data[32] = lut_32_ff;
    end
    else begin : no_ff_32
        assign out_data[32] = lut_32_out;
    end
    endgenerate
    
    
    
    // LUT : 33
    wire [15:0] lut_33_table = 16'b1101010001000000;
    wire [3:0] lut_33_select = {
                             in_data[135],
                             in_data[134],
                             in_data[133],
                             in_data[132]};
    
    wire lut_33_out = lut_33_table[lut_33_select];
    
    generate
    if ( USE_REG ) begin : ff_33
        reg   lut_33_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_33_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_33_ff <= lut_33_out;
            end
        end
        
        assign out_data[33] = lut_33_ff;
    end
    else begin : no_ff_33
        assign out_data[33] = lut_33_out;
    end
    endgenerate
    
    
    
    // LUT : 34
    wire [15:0] lut_34_table = 16'b1101010101000100;
    wire [3:0] lut_34_select = {
                             in_data[139],
                             in_data[138],
                             in_data[137],
                             in_data[136]};
    
    wire lut_34_out = lut_34_table[lut_34_select];
    
    generate
    if ( USE_REG ) begin : ff_34
        reg   lut_34_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_34_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_34_ff <= lut_34_out;
            end
        end
        
        assign out_data[34] = lut_34_ff;
    end
    else begin : no_ff_34
        assign out_data[34] = lut_34_out;
    end
    endgenerate
    
    
    
    // LUT : 35
    wire [15:0] lut_35_table = 16'b1000111100001110;
    wire [3:0] lut_35_select = {
                             in_data[143],
                             in_data[142],
                             in_data[141],
                             in_data[140]};
    
    wire lut_35_out = lut_35_table[lut_35_select];
    
    generate
    if ( USE_REG ) begin : ff_35
        reg   lut_35_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_35_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_35_ff <= lut_35_out;
            end
        end
        
        assign out_data[35] = lut_35_ff;
    end
    else begin : no_ff_35
        assign out_data[35] = lut_35_out;
    end
    endgenerate
    
    
    
    // LUT : 36
    wire [15:0] lut_36_table = 16'b0100110100000100;
    wire [3:0] lut_36_select = {
                             in_data[147],
                             in_data[146],
                             in_data[145],
                             in_data[144]};
    
    wire lut_36_out = lut_36_table[lut_36_select];
    
    generate
    if ( USE_REG ) begin : ff_36
        reg   lut_36_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_36_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_36_ff <= lut_36_out;
            end
        end
        
        assign out_data[36] = lut_36_ff;
    end
    else begin : no_ff_36
        assign out_data[36] = lut_36_out;
    end
    endgenerate
    
    
    
    // LUT : 37
    wire [15:0] lut_37_table = 16'b0101000101110011;
    wire [3:0] lut_37_select = {
                             in_data[151],
                             in_data[150],
                             in_data[149],
                             in_data[148]};
    
    wire lut_37_out = lut_37_table[lut_37_select];
    
    generate
    if ( USE_REG ) begin : ff_37
        reg   lut_37_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_37_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_37_ff <= lut_37_out;
            end
        end
        
        assign out_data[37] = lut_37_ff;
    end
    else begin : no_ff_37
        assign out_data[37] = lut_37_out;
    end
    endgenerate
    
    
    
    // LUT : 38
    wire [15:0] lut_38_table = 16'b0000101100111111;
    wire [3:0] lut_38_select = {
                             in_data[155],
                             in_data[154],
                             in_data[153],
                             in_data[152]};
    
    wire lut_38_out = lut_38_table[lut_38_select];
    
    generate
    if ( USE_REG ) begin : ff_38
        reg   lut_38_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_38_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_38_ff <= lut_38_out;
            end
        end
        
        assign out_data[38] = lut_38_ff;
    end
    else begin : no_ff_38
        assign out_data[38] = lut_38_out;
    end
    endgenerate
    
    
    
    // LUT : 39
    wire [15:0] lut_39_table = 16'b0000011100010111;
    wire [3:0] lut_39_select = {
                             in_data[159],
                             in_data[158],
                             in_data[157],
                             in_data[156]};
    
    wire lut_39_out = lut_39_table[lut_39_select];
    
    generate
    if ( USE_REG ) begin : ff_39
        reg   lut_39_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_39_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_39_ff <= lut_39_out;
            end
        end
        
        assign out_data[39] = lut_39_ff;
    end
    else begin : no_ff_39
        assign out_data[39] = lut_39_out;
    end
    endgenerate
    
    
endmodule



module MnistLutSimple_sub8
        #(
            parameter USER_WIDTH = 0,
            parameter USE_REG    = 1,
            parameter INIT_REG   = 1'bx,
            parameter DEVICE     = "RTL",
            
            parameter USER_BITS  = USER_WIDTH > 0 ? USER_WIDTH : 1
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [USER_BITS-1:0]  in_user,
            input  wire [         39:0]  in_data,
            input  wire                  in_valid,
            
            output wire [USER_BITS-1:0]  out_user,
            output wire [          9:0]  out_data,
            output wire                  out_valid
        );
    
    MnistLutSimple_sub8_base
            #(
                .USE_REG   (USE_REG),
                .INIT_REG  (INIT_REG),
                .DEVICE    (DEVICE)
            )
        i_MnistLutSimple_sub8_base
            (
                .reset     (reset),
                .clk       (clk),
                .cke       (cke),
                
                .in_data   (in_data),
                .out_data  (out_data)
            );
    
    generate
    if ( USE_REG ) begin : ff
        reg   [USER_BITS-1:0]  reg_out_user;
        reg                    reg_out_valid;
        always @(posedge clk) begin
            if ( reset ) begin
                reg_out_user  <= {USER_BITS{1'bx}};
                reg_out_valid <= 1'b0;
            end
            else if ( cke ) begin
                reg_out_user  <= in_user;
                reg_out_valid <= in_valid;
            end
        end
        assign out_user  = reg_out_user;
        assign out_valid = reg_out_valid;
    end
    else begin : no_ff
        assign out_user  = in_user;
        assign out_valid = in_valid;
    end
    endgenerate
    
    
endmodule




module MnistLutSimple_sub8_base
        #(
            parameter USE_REG  = 1,
            parameter INIT_REG = 1'bx,
            parameter DEVICE   = "RTL"
        )
        (
            input  wire         reset,
            input  wire         clk,
            input  wire         cke,
            
            input  wire [39:0]  in_data,
            output wire [9:0]  out_data
        );
    
    
    // LUT : 0
    wire [15:0] lut_0_table = 16'b1110100010000000;
    wire [3:0] lut_0_select = {
                             in_data[3],
                             in_data[2],
                             in_data[1],
                             in_data[0]};
    
    wire lut_0_out = lut_0_table[lut_0_select];
    
    generate
    if ( USE_REG ) begin : ff_0
        reg   lut_0_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_0_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_0_ff <= lut_0_out;
            end
        end
        
        assign out_data[0] = lut_0_ff;
    end
    else begin : no_ff_0
        assign out_data[0] = lut_0_out;
    end
    endgenerate
    
    
    
    // LUT : 1
    wire [15:0] lut_1_table = 16'b1110100010000000;
    wire [3:0] lut_1_select = {
                             in_data[7],
                             in_data[6],
                             in_data[5],
                             in_data[4]};
    
    wire lut_1_out = lut_1_table[lut_1_select];
    
    generate
    if ( USE_REG ) begin : ff_1
        reg   lut_1_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_1_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_1_ff <= lut_1_out;
            end
        end
        
        assign out_data[1] = lut_1_ff;
    end
    else begin : no_ff_1
        assign out_data[1] = lut_1_out;
    end
    endgenerate
    
    
    
    // LUT : 2
    wire [15:0] lut_2_table = 16'b1110100010000000;
    wire [3:0] lut_2_select = {
                             in_data[11],
                             in_data[10],
                             in_data[9],
                             in_data[8]};
    
    wire lut_2_out = lut_2_table[lut_2_select];
    
    generate
    if ( USE_REG ) begin : ff_2
        reg   lut_2_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_2_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_2_ff <= lut_2_out;
            end
        end
        
        assign out_data[2] = lut_2_ff;
    end
    else begin : no_ff_2
        assign out_data[2] = lut_2_out;
    end
    endgenerate
    
    
    
    // LUT : 3
    wire [15:0] lut_3_table = 16'b1110100010000000;
    wire [3:0] lut_3_select = {
                             in_data[15],
                             in_data[14],
                             in_data[13],
                             in_data[12]};
    
    wire lut_3_out = lut_3_table[lut_3_select];
    
    generate
    if ( USE_REG ) begin : ff_3
        reg   lut_3_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_3_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_3_ff <= lut_3_out;
            end
        end
        
        assign out_data[3] = lut_3_ff;
    end
    else begin : no_ff_3
        assign out_data[3] = lut_3_out;
    end
    endgenerate
    
    
    
    // LUT : 4
    wire [15:0] lut_4_table = 16'b1110100010000000;
    wire [3:0] lut_4_select = {
                             in_data[19],
                             in_data[18],
                             in_data[17],
                             in_data[16]};
    
    wire lut_4_out = lut_4_table[lut_4_select];
    
    generate
    if ( USE_REG ) begin : ff_4
        reg   lut_4_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_4_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_4_ff <= lut_4_out;
            end
        end
        
        assign out_data[4] = lut_4_ff;
    end
    else begin : no_ff_4
        assign out_data[4] = lut_4_out;
    end
    endgenerate
    
    
    
    // LUT : 5
    wire [15:0] lut_5_table = 16'b1110100010000000;
    wire [3:0] lut_5_select = {
                             in_data[23],
                             in_data[22],
                             in_data[21],
                             in_data[20]};
    
    wire lut_5_out = lut_5_table[lut_5_select];
    
    generate
    if ( USE_REG ) begin : ff_5
        reg   lut_5_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_5_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_5_ff <= lut_5_out;
            end
        end
        
        assign out_data[5] = lut_5_ff;
    end
    else begin : no_ff_5
        assign out_data[5] = lut_5_out;
    end
    endgenerate
    
    
    
    // LUT : 6
    wire [15:0] lut_6_table = 16'b1110100010000000;
    wire [3:0] lut_6_select = {
                             in_data[27],
                             in_data[26],
                             in_data[25],
                             in_data[24]};
    
    wire lut_6_out = lut_6_table[lut_6_select];
    
    generate
    if ( USE_REG ) begin : ff_6
        reg   lut_6_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_6_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_6_ff <= lut_6_out;
            end
        end
        
        assign out_data[6] = lut_6_ff;
    end
    else begin : no_ff_6
        assign out_data[6] = lut_6_out;
    end
    endgenerate
    
    
    
    // LUT : 7
    wire [15:0] lut_7_table = 16'b1110100010000000;
    wire [3:0] lut_7_select = {
                             in_data[31],
                             in_data[30],
                             in_data[29],
                             in_data[28]};
    
    wire lut_7_out = lut_7_table[lut_7_select];
    
    generate
    if ( USE_REG ) begin : ff_7
        reg   lut_7_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_7_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_7_ff <= lut_7_out;
            end
        end
        
        assign out_data[7] = lut_7_ff;
    end
    else begin : no_ff_7
        assign out_data[7] = lut_7_out;
    end
    endgenerate
    
    
    
    // LUT : 8
    wire [15:0] lut_8_table = 16'b1110100010000000;
    wire [3:0] lut_8_select = {
                             in_data[35],
                             in_data[34],
                             in_data[33],
                             in_data[32]};
    
    wire lut_8_out = lut_8_table[lut_8_select];
    
    generate
    if ( USE_REG ) begin : ff_8
        reg   lut_8_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_8_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_8_ff <= lut_8_out;
            end
        end
        
        assign out_data[8] = lut_8_ff;
    end
    else begin : no_ff_8
        assign out_data[8] = lut_8_out;
    end
    endgenerate
    
    
    
    // LUT : 9
    wire [15:0] lut_9_table = 16'b1110100010000000;
    wire [3:0] lut_9_select = {
                             in_data[39],
                             in_data[38],
                             in_data[37],
                             in_data[36]};
    
    wire lut_9_out = lut_9_table[lut_9_select];
    
    generate
    if ( USE_REG ) begin : ff_9
        reg   lut_9_ff;
        always @(posedge clk) begin
            if ( reset ) begin
                lut_9_ff <= INIT_REG;
            end
            else if ( cke ) begin
                lut_9_ff <= lut_9_out;
            end
        end
        
        assign out_data[9] = lut_9_ff;
    end
    else begin : no_ff_9
        assign out_data[9] = lut_9_out;
    end
    endgenerate
    
    
endmodule

